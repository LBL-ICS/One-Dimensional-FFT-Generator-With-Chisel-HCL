module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 72:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[Arithmetic.scala 72:34]
  wire [8:0] result = _result_T_2[8:0]; // @[Arithmetic.scala 71:22 72:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 73:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 74:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 8'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module full_adder(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [24:0] result = _result_T_1[24:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[23:0]; // @[Arithmetic.scala 59:23]
  assign io_out_c = result[24]; // @[Arithmetic.scala 60:23]
endmodule
module twoscomplement_1(
  input  [23:0] io_in,
  output [23:0] io_out
);
  wire [23:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 24'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module shifter(
  input  [23:0] io_in_a,
  input  [4:0]  io_in_b,
  output [23:0] io_out_s
);
  wire [23:0] _result_T = io_in_a >> io_in_b; // @[Arithmetic.scala 42:25]
  wire [54:0] _GEN_0 = {{31'd0}, _result_T}; // @[Arithmetic.scala 41:26 42:14 44:14]
  assign io_out_s = _GEN_0[23:0]; // @[Arithmetic.scala 39:22]
endmodule
module leadingOneDetector(
  input  [23:0] io_in,
  output [4:0]  io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  assign io_out = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
endmodule
module FP_adder(
  input         clock,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 76:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 76:24]
  wire [7:0] complement_io_in; // @[FPArithmetic.scala 82:28]
  wire [7:0] complement_io_out; // @[FPArithmetic.scala 82:28]
  wire [23:0] adder_io_in_a; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_in_b; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_out_s; // @[FPArithmetic.scala 86:23]
  wire  adder_io_out_c; // @[FPArithmetic.scala 86:23]
  wire [23:0] complementN_0_io_in; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_0_io_out; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_1_io_in; // @[FPArithmetic.scala 94:31]
  wire [23:0] complementN_1_io_out; // @[FPArithmetic.scala 94:31]
  wire [23:0] shifter_io_in_a; // @[FPArithmetic.scala 98:25]
  wire [4:0] shifter_io_in_b; // @[FPArithmetic.scala 98:25]
  wire [23:0] shifter_io_out_s; // @[FPArithmetic.scala 98:25]
  wire [23:0] complementN_2_io_in; // @[FPArithmetic.scala 143:31]
  wire [23:0] complementN_2_io_out; // @[FPArithmetic.scala 143:31]
  wire [23:0] leadingOneFinder_io_in; // @[FPArithmetic.scala 163:34]
  wire [4:0] leadingOneFinder_io_out; // @[FPArithmetic.scala 163:34]
  wire [7:0] subber2_io_in_a; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_in_b; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_out_s; // @[FPArithmetic.scala 165:25]
  wire  subber2_io_out_c; // @[FPArithmetic.scala 165:25]
  wire  sign_0 = io_in_a[31]; // @[FPArithmetic.scala 38:23]
  wire  sign_1 = io_in_b[31]; // @[FPArithmetic.scala 39:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 43:62]
  wire [8:0] _GEN_31 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:34]
  wire [8:0] _GEN_0 = _GEN_31 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:68 44:14 46:14]
  wire [8:0] _GEN_32 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:34]
  wire [8:0] _GEN_1 = _GEN_32 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:68 49:14 51:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 56:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 57:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FPArithmetic.scala 61:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FPArithmetic.scala 62:26]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] out_exp = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  wire [7:0] sub_exp = subber_io_out_c ? complement_io_out : subber_io_out_s; // @[FPArithmetic.scala 104:34 106:15 116:15]
  wire  out_s = subber_io_out_c ? sign_1 : sign_0; // @[FPArithmetic.scala 104:34 107:13 117:13]
  wire [22:0] out_frac = subber_io_out_c ? frac_1 : frac_0; // @[FPArithmetic.scala 104:34 108:16 118:16]
  wire [23:0] _GEN_8 = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  wire [23:0] _GEN_9 = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  wire  _new_s_T = ~adder_io_out_c; // @[FPArithmetic.scala 138:15]
  wire  _D_T_1 = sign_0 ^ sign_1; // @[FPArithmetic.scala 151:39]
  wire  D = _new_s_T | sign_0 ^ sign_1; // @[FPArithmetic.scala 151:28]
  wire  E = _new_s_T & ~adder_io_out_s[23] | _new_s_T & ~_D_T_1 | adder_io_out_c & adder_io_out_s[23] & _D_T_1; // @[FPArithmetic.scala 154:99]
  wire  _GEN_25 = sub_exp >= 8'h17 ? out_s : ~adder_io_out_c & sign_0 | sign_0 & sign_1 | ~adder_io_out_c & sign_1; // @[FPArithmetic.scala 138:11 173:39 174:13]
  wire  new_s = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 1'h0 : _GEN_25; // @[FPArithmetic.scala 169:62 170:13]
  wire [23:0] adder_result = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  wire [4:0] _subber2_io_in_b_T_1 = 5'h18 - leadingOneFinder_io_out; // @[FPArithmetic.scala 167:42]
  wire [8:0] _GEN_33 = {{1'd0}, out_exp}; // @[FPArithmetic.scala 181:20]
  wire [23:0] _new_out_frac_T_2 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 183:51]
  wire [7:0] _new_out_exp_T_3 = out_exp + 8'h1; // @[FPArithmetic.scala 185:32]
  wire [8:0] _GEN_13 = _GEN_33 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_T_3}; // @[FPArithmetic.scala 181:56 182:21 185:21]
  wire [23:0] _GEN_14 = _GEN_33 == _T_2 ? _new_out_frac_T_2 : {{1'd0}, adder_result[23:1]}; // @[FPArithmetic.scala 181:56 183:22 186:22]
  wire [53:0] _GEN_2 = {{31'd0}, adder_result[22:0]}; // @[FPArithmetic.scala 197:57]
  wire [53:0] _new_out_frac_T_7 = _GEN_2 << _subber2_io_in_b_T_1; // @[FPArithmetic.scala 197:57]
  wire [7:0] _GEN_15 = subber2_io_out_c ? 8'h1 : subber2_io_out_s; // @[FPArithmetic.scala 192:39 193:23 196:23]
  wire [53:0] _GEN_16 = subber2_io_out_c ? 54'h400000 : _new_out_frac_T_7; // @[FPArithmetic.scala 192:39 194:24 197:24]
  wire [7:0] _GEN_17 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:0
    ]) ? 8'h0 : _GEN_15; // @[FPArithmetic.scala 189:141 190:21]
  wire [53:0] _GEN_18 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:
    0]) ? 54'h0 : _GEN_16; // @[FPArithmetic.scala 189:141 139:18]
  wire [7:0] _GEN_19 = D ? _GEN_17 : 8'h0; // @[FPArithmetic.scala 140:17 188:26]
  wire [53:0] _GEN_20 = D ? _GEN_18 : 54'h0; // @[FPArithmetic.scala 139:18 188:26]
  wire [8:0] _GEN_21 = ~D ? _GEN_13 : {{1'd0}, _GEN_19}; // @[FPArithmetic.scala 180:26]
  wire [53:0] _GEN_22 = ~D ? {{30'd0}, _GEN_14} : _GEN_20; // @[FPArithmetic.scala 180:26]
  wire [8:0] _GEN_23 = E ? {{1'd0}, out_exp} : _GEN_21; // @[FPArithmetic.scala 177:26 178:19]
  wire [53:0] _GEN_24 = E ? {{31'd0}, adder_result[22:0]} : _GEN_22; // @[FPArithmetic.scala 177:26 179:20]
  wire [53:0] _GEN_26 = sub_exp >= 8'h17 ? {{31'd0}, out_frac} : _GEN_24; // @[FPArithmetic.scala 173:39 175:20]
  wire [8:0] _GEN_27 = sub_exp >= 8'h17 ? {{1'd0}, out_exp} : _GEN_23; // @[FPArithmetic.scala 173:39 176:19]
  wire [8:0] _GEN_29 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 9'h0 : _GEN_27; // @[FPArithmetic.scala 169:62 171:19]
  wire [53:0] _GEN_30 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 54'h0 : _GEN_26; // @[FPArithmetic.scala 169:62 172:20]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 201:24]
  wire [7:0] new_out_exp = _GEN_29[7:0]; // @[FPArithmetic.scala 137:27]
  wire [8:0] _reg_out_s_T = {new_s,new_out_exp}; // @[FPArithmetic.scala 202:24]
  wire [22:0] new_out_frac = _GEN_30[22:0]; // @[FPArithmetic.scala 136:28]
  full_subber subber ( // @[FPArithmetic.scala 76:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complement ( // @[FPArithmetic.scala 82:28]
    .io_in(complement_io_in),
    .io_out(complement_io_out)
  );
  full_adder adder ( // @[FPArithmetic.scala 86:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  twoscomplement_1 complementN_0 ( // @[FPArithmetic.scala 92:31]
    .io_in(complementN_0_io_in),
    .io_out(complementN_0_io_out)
  );
  twoscomplement_1 complementN_1 ( // @[FPArithmetic.scala 94:31]
    .io_in(complementN_1_io_in),
    .io_out(complementN_1_io_out)
  );
  shifter shifter ( // @[FPArithmetic.scala 98:25]
    .io_in_a(shifter_io_in_a),
    .io_in_b(shifter_io_in_b),
    .io_out_s(shifter_io_out_s)
  );
  twoscomplement_1 complementN_2 ( // @[FPArithmetic.scala 143:31]
    .io_in(complementN_2_io_in),
    .io_out(complementN_2_io_out)
  );
  leadingOneDetector leadingOneFinder ( // @[FPArithmetic.scala 163:34]
    .io_in(leadingOneFinder_io_in),
    .io_out(leadingOneFinder_io_out)
  );
  full_subber subber2 ( // @[FPArithmetic.scala 165:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 204:14]
  assign subber_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  assign complement_io_in = subber_io_out_s; // @[FPArithmetic.scala 83:22]
  assign adder_io_in_a = sign_0 & ~sign_1 ? complementN_0_io_out : _GEN_8; // @[FPArithmetic.scala 127:45 128:21]
  assign adder_io_in_b = sign_1 & ~sign_0 ? complementN_1_io_out : _GEN_9; // @[FPArithmetic.scala 131:45 132:21]
  assign complementN_0_io_in = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  assign complementN_1_io_in = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  assign shifter_io_in_a = subber_io_out_c ? whole_frac_0 : whole_frac_1; // @[FPArithmetic.scala 104:34 109:23 119:23]
  assign shifter_io_in_b = sub_exp[4:0];
  assign complementN_2_io_in = adder_io_out_s; // @[FPArithmetic.scala 144:25]
  assign leadingOneFinder_io_in = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  assign subber2_io_in_a = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  assign subber2_io_in_b = {{3'd0}, _subber2_io_in_b_T_1}; // @[FPArithmetic.scala 167:21]
  always @(posedge clock) begin
    reg_out_s <= {_reg_out_s_T,new_out_frac}; // @[FPArithmetic.scala 202:39]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexAdder(
  input         clock,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_adder_clock; // @[FPComplex.scala 20:25]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 20:25]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 20:25]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 20:25]
  wire  FP_adder_1_clock; // @[FPComplex.scala 20:25]
  wire [31:0] FP_adder_1_io_in_a; // @[FPComplex.scala 20:25]
  wire [31:0] FP_adder_1_io_in_b; // @[FPComplex.scala 20:25]
  wire [31:0] FP_adder_1_io_out_s; // @[FPComplex.scala 20:25]
  FP_adder FP_adder ( // @[FPComplex.scala 20:25]
    .clock(FP_adder_clock),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_adder FP_adder_1 ( // @[FPComplex.scala 20:25]
    .clock(FP_adder_1_clock),
    .io_in_a(FP_adder_1_io_in_a),
    .io_in_b(FP_adder_1_io_in_b),
    .io_out_s(FP_adder_1_io_out_s)
  );
  assign io_out_s_Re = FP_adder_io_out_s; // @[FPComplex.scala 27:17]
  assign io_out_s_Im = FP_adder_1_io_out_s; // @[FPComplex.scala 28:17]
  assign FP_adder_clock = clock;
  assign FP_adder_io_in_a = io_in_a_Re; // @[FPComplex.scala 23:23]
  assign FP_adder_io_in_b = io_in_b_Re; // @[FPComplex.scala 24:23]
  assign FP_adder_1_clock = clock;
  assign FP_adder_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 25:23]
  assign FP_adder_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 26:23]
endmodule
module FPComplexMultiAdder(
  input         clock,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  FPComplexAdder_clock; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 178:28]
  wire  FPComplexAdder_1_clock; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_1_io_in_a_Re; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_1_io_in_a_Im; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_1_io_in_b_Re; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_1_io_in_b_Im; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_1_io_out_s_Re; // @[FPComplex.scala 178:28]
  wire [31:0] FPComplexAdder_1_io_out_s_Im; // @[FPComplex.scala 178:28]
  FPComplexAdder FPComplexAdder ( // @[FPComplex.scala 178:28]
    .clock(FPComplexAdder_clock),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_1 ( // @[FPComplex.scala 178:28]
    .clock(FPComplexAdder_1_clock),
    .io_in_a_Re(FPComplexAdder_1_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_1_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_1_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_1_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_1_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_1_io_out_s_Im)
  );
  assign io_out_Re = FPComplexAdder_1_io_out_s_Re; // @[FPComplex.scala 233:12]
  assign io_out_Im = FPComplexAdder_1_io_out_s_Im; // @[FPComplex.scala 233:12]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_io_in_a_Re = io_in_0_Re; // @[FPComplex.scala 195:38]
  assign FPComplexAdder_io_in_a_Im = io_in_0_Im; // @[FPComplex.scala 195:38]
  assign FPComplexAdder_io_in_b_Re = io_in_1_Re; // @[FPComplex.scala 196:38]
  assign FPComplexAdder_io_in_b_Im = io_in_1_Im; // @[FPComplex.scala 196:38]
  assign FPComplexAdder_1_clock = clock;
  assign FPComplexAdder_1_io_in_a_Re = FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 205:40]
  assign FPComplexAdder_1_io_in_a_Im = FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 205:40]
  assign FPComplexAdder_1_io_in_b_Re = io_in_2_Re; // @[FPComplex.scala 190:39]
  assign FPComplexAdder_1_io_in_b_Im = io_in_2_Im; // @[FPComplex.scala 190:39]
endmodule
module FP_subber(
  input         clock,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FPArithmetic.scala 216:26]
  wire [31:0] FP_adder_io_in_a; // @[FPArithmetic.scala 216:26]
  wire [31:0] FP_adder_io_in_b; // @[FPArithmetic.scala 216:26]
  wire [31:0] FP_adder_io_out_s; // @[FPArithmetic.scala 216:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FPArithmetic.scala 219:23]
  FP_adder FP_adder ( // @[FPArithmetic.scala 216:26]
    .clock(FP_adder_clock),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FPArithmetic.scala 222:14]
  assign FP_adder_clock = clock;
  assign FP_adder_io_in_a = io_in_a; // @[FPArithmetic.scala 220:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FPArithmetic.scala 219:39]
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[Arithmetic.scala 84:23]
endmodule
module full_adder_14(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [8:0] result = _result_T_1[8:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 59:23]
endmodule
module FP_multiplier(
  input         clock,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FPArithmetic.scala 290:28]
  wire [23:0] multiplier_io_in_b; // @[FPArithmetic.scala 290:28]
  wire [47:0] multiplier_io_out_s; // @[FPArithmetic.scala 290:28]
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 295:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 295:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 295:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 295:24]
  wire [7:0] complementN_io_in; // @[FPArithmetic.scala 301:29]
  wire [7:0] complementN_io_out; // @[FPArithmetic.scala 301:29]
  wire [7:0] adderN_io_in_a; // @[FPArithmetic.scala 305:24]
  wire [7:0] adderN_io_in_b; // @[FPArithmetic.scala 305:24]
  wire [7:0] adderN_io_out_s; // @[FPArithmetic.scala 305:24]
  wire  s_0 = io_in_a[31]; // @[FPArithmetic.scala 255:20]
  wire  s_1 = io_in_b[31]; // @[FPArithmetic.scala 256:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 260:62]
  wire [8:0] _GEN_13 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 260:34]
  wire [8:0] _GEN_0 = _GEN_13 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 260:68 261:14 263:14]
  wire [8:0] _GEN_14 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 265:34]
  wire [8:0] _GEN_1 = _GEN_14 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 265:68 266:14 268:14]
  wire [22:0] exp_check_0 = {{15'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 271:25 272:18]
  wire [22:0] _cond_holder_T_1 = exp_check_0 + 23'h1; // @[FPArithmetic.scala 276:34]
  wire [22:0] exp_check_1 = {{15'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 271:25 273:18]
  wire [22:0] _cond_holder_T_3 = 23'h7f - exp_check_1; // @[FPArithmetic.scala 276:80]
  wire [22:0] _cond_holder_T_4 = ~_cond_holder_T_3; // @[FPArithmetic.scala 276:42]
  wire [22:0] _cond_holder_T_6 = _cond_holder_T_1 + _cond_holder_T_4; // @[FPArithmetic.scala 276:40]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 280:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 281:23]
  wire  new_s = s_0 ^ s_1; // @[FPArithmetic.scala 312:19]
  wire [7:0] _new_exp_T_1 = adderN_io_out_s + 8'h1; // @[FPArithmetic.scala 323:34]
  wire [22:0] _cond_holder_T_8 = exp_check_0 + 23'h2; // @[FPArithmetic.scala 325:36]
  wire [22:0] _cond_holder_T_13 = _cond_holder_T_8 + _cond_holder_T_4; // @[FPArithmetic.scala 325:42]
  wire [23:0] _new_mant_T_2 = {multiplier_io_out_s[46:24], 1'h0}; // @[FPArithmetic.scala 331:73]
  wire [7:0] _GEN_2 = multiplier_io_out_s[47] ? _new_exp_T_1 : adderN_io_out_s; // @[FPArithmetic.scala 322:60 323:15 328:15]
  wire [22:0] cond_holder = multiplier_io_out_s[47] ? _cond_holder_T_13 : _cond_holder_T_6; // @[FPArithmetic.scala 322:60 325:19 330:19]
  wire [23:0] _GEN_5 = multiplier_io_out_s[47] ? {{1'd0}, multiplier_io_out_s[46:24]} : _new_mant_T_2; // @[FPArithmetic.scala 322:60 326:16 331:16]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 333:24]
  wire [22:0] _T_12 = ~cond_holder; // @[FPArithmetic.scala 334:51]
  wire [22:0] _T_14 = 23'h1 + _T_12; // @[FPArithmetic.scala 334:49]
  wire [22:0] _GEN_15 = {{14'd0}, _T_2}; // @[FPArithmetic.scala 334:42]
  wire [8:0] _GEN_6 = cond_holder > _GEN_15 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 339:61 340:15]
  wire [8:0] _GEN_9 = _GEN_15 >= _T_14 ? 9'h1 : _GEN_6; // @[FPArithmetic.scala 334:67 335:15]
  wire [7:0] new_exp = _GEN_9[7:0]; // @[FPArithmetic.scala 315:23]
  wire [23:0] _new_mant_T_4 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 341:45]
  wire [23:0] _GEN_7 = cond_holder > _GEN_15 ? _new_mant_T_4 : _GEN_5; // @[FPArithmetic.scala 339:61 341:16]
  wire [23:0] _GEN_10 = _GEN_15 >= _T_14 ? 24'h400000 : _GEN_7; // @[FPArithmetic.scala 334:67 336:16]
  wire [22:0] new_mant = _GEN_10[22:0]; // @[FPArithmetic.scala 317:24]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_exp,new_mant}; // @[FPArithmetic.scala 337:37]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 259:19]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 259:19]
  multiplier multiplier ( // @[FPArithmetic.scala 290:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FPArithmetic.scala 295:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FPArithmetic.scala 301:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder_14 adderN ( // @[FPArithmetic.scala 305:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 349:14]
  assign multiplier_io_in_a = {1'h1,frac_0}; // @[FPArithmetic.scala 285:24]
  assign multiplier_io_in_b = {1'h1,frac_1}; // @[FPArithmetic.scala 286:24]
  assign subber_io_in_a = 8'h7f; // @[FPArithmetic.scala 296:20]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 259:19]
  assign complementN_io_in = subber_io_out_s; // @[FPArithmetic.scala 302:23]
  assign adderN_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 259:19]
  assign adderN_io_in_b = complementN_io_out; // @[FPArithmetic.scala 307:20]
  always @(posedge clock) begin
    if (exp_0 == 8'h0 | exp_1 == 8'h0) begin // @[FPArithmetic.scala 344:43]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 345:17]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 347:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult_reducable(
  input         clock,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FP_subber_clock; // @[FPComplex.scala 84:24]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 84:24]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 84:24]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 84:24]
  wire  FP_adder_clock; // @[FPComplex.scala 85:24]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 85:24]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 85:24]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 85:24]
  wire  FP_multiplier_clock; // @[FPComplex.scala 155:28]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 155:28]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 155:28]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 155:28]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 155:28]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 155:28]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 155:28]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 155:28]
  wire  sign_0 = io_in_a_Re[31]; // @[FPComplex.scala 87:26]
  wire  sign_1 = io_in_a_Im[31]; // @[FPComplex.scala 88:26]
  wire [7:0] exp_0 = io_in_a_Re[30:23]; // @[FPComplex.scala 90:25]
  wire [7:0] exp_1 = io_in_a_Im[30:23]; // @[FPComplex.scala 91:25]
  wire [22:0] frac_0 = io_in_a_Re[22:0]; // @[FPComplex.scala 93:26]
  wire [22:0] frac_1 = io_in_a_Im[22:0]; // @[FPComplex.scala 94:26]
  wire [7:0] _new_exp1_0_T_1 = exp_0 - 8'h1; // @[FPComplex.scala 103:31]
  wire [7:0] new_exp1_0 = exp_0 != 8'h0 ? _new_exp1_0_T_1 : exp_0; // @[FPComplex.scala 102:27 103:21 105:21]
  wire [7:0] _new_exp1_1_T_1 = exp_1 - 8'h1; // @[FPComplex.scala 108:31]
  wire [7:0] new_exp1_1 = exp_1 != 8'h0 ? _new_exp1_1_T_1 : exp_1; // @[FPComplex.scala 107:27 108:21 110:21]
  reg [31:0] regs1_0; // @[FPComplex.scala 130:22]
  reg [31:0] regs1_1; // @[FPComplex.scala 130:22]
  wire [8:0] _regs1_0_T = {sign_0,new_exp1_0}; // @[FPComplex.scala 131:27]
  wire [8:0] _regs1_1_T = {sign_1,new_exp1_1}; // @[FPComplex.scala 132:27]
  FP_subber FP_subber ( // @[FPComplex.scala 84:24]
    .clock(FP_subber_clock),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 85:24]
    .clock(FP_adder_clock),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 155:28]
    .clock(FP_multiplier_clock),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 155:28]
    .clock(FP_multiplier_1_clock),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 169:17]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 170:17]
  assign FP_subber_clock = clock;
  assign FP_subber_io_in_a = regs1_0; // @[FPComplex.scala 128:28 133:23]
  assign FP_subber_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 128:28 163:23]
  assign FP_adder_clock = clock;
  assign FP_adder_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 128:28 162:23]
  assign FP_adder_io_in_b = regs1_1; // @[FPComplex.scala 128:28 134:23]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 158:31]
  assign FP_multiplier_io_in_b = io_in_b_Im; // @[FPComplex.scala 159:31]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 160:31]
  assign FP_multiplier_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 161:31]
  always @(posedge clock) begin
    regs1_0 <= {_regs1_0_T,frac_0}; // @[FPComplex.scala 131:42]
    regs1_1 <= {_regs1_1_T,frac_1}; // @[FPComplex.scala 132:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs1_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs1_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DFT_r_V1(
  input         clock,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexMultiAdder_clock; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_in_2_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_in_2_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 430:26]
  wire  FPComplexMultiAdder_1_clock; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_2_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_2_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 430:26]
  wire  FPComplexMultiAdder_2_clock; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_in_1_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_in_1_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_in_2_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_in_2_Im; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 430:26]
  wire [31:0] FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 430:26]
  wire  FPComplexMult_reducable_clock; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_io_in_a_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_io_in_a_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_io_in_b_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_io_out_s_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_io_out_s_Im; // @[FFTDesigns.scala 435:28]
  wire  FPComplexMult_reducable_1_clock; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_a_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_a_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_b_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_1_io_out_s_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_1_io_out_s_Im; // @[FFTDesigns.scala 435:28]
  wire  FPComplexMult_reducable_2_clock; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_a_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_a_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_b_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_2_io_out_s_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_2_io_out_s_Im; // @[FFTDesigns.scala 435:28]
  wire  FPComplexMult_reducable_3_clock; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_a_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_a_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_b_Im; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_3_io_out_s_Re; // @[FFTDesigns.scala 435:28]
  wire [31:0] FPComplexMult_reducable_3_io_out_s_Im; // @[FFTDesigns.scala 435:28]
  reg [31:0] reg_syncs_0_0_Re; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_0_0_Im; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_0_1_Re; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_0_1_Im; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_0_2_Re; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_0_2_Im; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_1_0_Re; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_1_0_Im; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_1_1_Re; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_1_1_Im; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_1_2_Re; // @[FFTDesigns.scala 445:23]
  reg [31:0] reg_syncs_1_2_Im; // @[FFTDesigns.scala 445:23]
  FPComplexMultiAdder FPComplexMultiAdder ( // @[FFTDesigns.scala 430:26]
    .clock(FPComplexMultiAdder_clock),
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_io_in_1_Im),
    .io_in_2_Re(FPComplexMultiAdder_io_in_2_Re),
    .io_in_2_Im(FPComplexMultiAdder_io_in_2_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 430:26]
    .clock(FPComplexMultiAdder_1_clock),
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_1_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_1_io_in_1_Im),
    .io_in_2_Re(FPComplexMultiAdder_1_io_in_2_Re),
    .io_in_2_Im(FPComplexMultiAdder_1_io_in_2_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder_2 ( // @[FFTDesigns.scala 430:26]
    .clock(FPComplexMultiAdder_2_clock),
    .io_in_0_Re(FPComplexMultiAdder_2_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_2_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_2_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_2_io_in_1_Im),
    .io_in_2_Re(FPComplexMultiAdder_2_io_in_2_Re),
    .io_in_2_Im(FPComplexMultiAdder_2_io_in_2_Im),
    .io_out_Re(FPComplexMultiAdder_2_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_2_io_out_Im)
  );
  FPComplexMult_reducable FPComplexMult_reducable ( // @[FFTDesigns.scala 435:28]
    .clock(FPComplexMult_reducable_clock),
    .io_in_a_Re(FPComplexMult_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_io_in_a_Im),
    .io_in_b_Im(FPComplexMult_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_io_out_s_Im)
  );
  FPComplexMult_reducable FPComplexMult_reducable_1 ( // @[FFTDesigns.scala 435:28]
    .clock(FPComplexMult_reducable_1_clock),
    .io_in_a_Re(FPComplexMult_reducable_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_1_io_in_a_Im),
    .io_in_b_Im(FPComplexMult_reducable_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_1_io_out_s_Im)
  );
  FPComplexMult_reducable FPComplexMult_reducable_2 ( // @[FFTDesigns.scala 435:28]
    .clock(FPComplexMult_reducable_2_clock),
    .io_in_a_Re(FPComplexMult_reducable_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_2_io_in_a_Im),
    .io_in_b_Im(FPComplexMult_reducable_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_2_io_out_s_Im)
  );
  FPComplexMult_reducable FPComplexMult_reducable_3 ( // @[FFTDesigns.scala 435:28]
    .clock(FPComplexMult_reducable_3_clock),
    .io_in_a_Re(FPComplexMult_reducable_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_3_io_in_a_Im),
    .io_in_b_Im(FPComplexMult_reducable_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_3_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 494:22 496:17]
  assign io_out_0_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 494:22 496:17]
  assign io_out_1_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 494:22 496:17]
  assign io_out_1_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 494:22 496:17]
  assign io_out_2_Re = FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 494:22 496:17]
  assign io_out_2_Im = FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 494:22 496:17]
  assign FPComplexMultiAdder_clock = clock;
  assign FPComplexMultiAdder_io_in_0_Re = reg_syncs_1_0_Re; // @[FFTDesigns.scala 460:30 462:28]
  assign FPComplexMultiAdder_io_in_0_Im = reg_syncs_1_0_Im; // @[FFTDesigns.scala 460:30 462:28]
  assign FPComplexMultiAdder_io_in_1_Re = reg_syncs_1_1_Re; // @[FFTDesigns.scala 460:30 462:28]
  assign FPComplexMultiAdder_io_in_1_Im = reg_syncs_1_1_Im; // @[FFTDesigns.scala 460:30 462:28]
  assign FPComplexMultiAdder_io_in_2_Re = reg_syncs_1_2_Re; // @[FFTDesigns.scala 460:30 462:28]
  assign FPComplexMultiAdder_io_in_2_Im = reg_syncs_1_2_Im; // @[FFTDesigns.scala 460:30 462:28]
  assign FPComplexMultiAdder_1_clock = clock;
  assign FPComplexMultiAdder_1_io_in_0_Re = reg_syncs_1_0_Re; // @[FFTDesigns.scala 460:30 464:30]
  assign FPComplexMultiAdder_1_io_in_0_Im = reg_syncs_1_0_Im; // @[FFTDesigns.scala 460:30 464:30]
  assign FPComplexMultiAdder_1_io_in_1_Re = FPComplexMult_reducable_io_out_s_Re; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_1_io_in_1_Im = FPComplexMult_reducable_io_out_s_Im; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_1_io_in_2_Re = FPComplexMult_reducable_1_io_out_s_Re; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_1_io_in_2_Im = FPComplexMult_reducable_1_io_out_s_Im; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_2_clock = clock;
  assign FPComplexMultiAdder_2_io_in_0_Re = reg_syncs_1_0_Re; // @[FFTDesigns.scala 460:30 464:30]
  assign FPComplexMultiAdder_2_io_in_0_Im = reg_syncs_1_0_Im; // @[FFTDesigns.scala 460:30 464:30]
  assign FPComplexMultiAdder_2_io_in_1_Re = FPComplexMult_reducable_2_io_out_s_Re; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_2_io_in_1_Im = FPComplexMult_reducable_2_io_out_s_Im; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_2_io_in_2_Re = FPComplexMult_reducable_3_io_out_s_Re; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMultiAdder_2_io_in_2_Im = FPComplexMult_reducable_3_io_out_s_Im; // @[FFTDesigns.scala 460:30 470:52]
  assign FPComplexMult_reducable_clock = clock;
  assign FPComplexMult_reducable_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_io_in_b_Im = 32'hbf5db3d6; // @[FFTDesigns.scala 441:29]
  assign FPComplexMult_reducable_1_clock = clock;
  assign FPComplexMult_reducable_1_io_in_a_Re = io_in_2_Re; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_1_io_in_a_Im = io_in_2_Im; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_1_io_in_b_Im = 32'h3f5db3d6; // @[FFTDesigns.scala 441:29]
  assign FPComplexMult_reducable_2_clock = clock;
  assign FPComplexMult_reducable_2_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_2_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_2_io_in_b_Im = 32'h3f5db3d6; // @[FFTDesigns.scala 441:29]
  assign FPComplexMult_reducable_3_clock = clock;
  assign FPComplexMult_reducable_3_io_in_a_Re = io_in_2_Re; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_3_io_in_a_Im = io_in_2_Im; // @[FFTDesigns.scala 409:24 418:33]
  assign FPComplexMult_reducable_3_io_in_b_Im = 32'hbf5db3d6; // @[FFTDesigns.scala 441:29]
  always @(posedge clock) begin
    reg_syncs_0_0_Re <= io_in_0_Re; // @[FFTDesigns.scala 451:29]
    reg_syncs_0_0_Im <= io_in_0_Im; // @[FFTDesigns.scala 451:29]
    reg_syncs_0_1_Re <= io_in_1_Re; // @[FFTDesigns.scala 451:29]
    reg_syncs_0_1_Im <= io_in_1_Im; // @[FFTDesigns.scala 451:29]
    reg_syncs_0_2_Re <= io_in_2_Re; // @[FFTDesigns.scala 451:29]
    reg_syncs_0_2_Im <= io_in_2_Im; // @[FFTDesigns.scala 451:29]
    reg_syncs_1_0_Re <= reg_syncs_0_0_Re; // @[FFTDesigns.scala 457:24]
    reg_syncs_1_0_Im <= reg_syncs_0_0_Im; // @[FFTDesigns.scala 457:24]
    reg_syncs_1_1_Re <= reg_syncs_0_1_Re; // @[FFTDesigns.scala 457:24]
    reg_syncs_1_1_Im <= reg_syncs_0_1_Im; // @[FFTDesigns.scala 457:24]
    reg_syncs_1_2_Re <= reg_syncs_0_2_Re; // @[FFTDesigns.scala 457:24]
    reg_syncs_1_2_Im <= reg_syncs_0_2_Im; // @[FFTDesigns.scala 457:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_syncs_0_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_syncs_0_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_syncs_0_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_syncs_0_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_syncs_0_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_syncs_0_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_syncs_1_0_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_syncs_1_0_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_syncs_1_1_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_syncs_1_1_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_syncs_1_2_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_syncs_1_2_Im = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationsBasic(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_1_Re = io_in_9_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_1_Im = io_in_9_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_2_Re = io_in_18_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_2_Im = io_in_18_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_3_Re = io_in_3_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_3_Im = io_in_3_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_4_Re = io_in_12_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_4_Im = io_in_12_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_5_Re = io_in_21_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_5_Im = io_in_21_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_6_Re = io_in_6_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_6_Im = io_in_6_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_7_Re = io_in_15_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_7_Im = io_in_15_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_8_Re = io_in_24_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_8_Im = io_in_24_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_9_Re = io_in_1_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_9_Im = io_in_1_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_10_Re = io_in_10_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_10_Im = io_in_10_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_11_Re = io_in_19_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_11_Im = io_in_19_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_12_Re = io_in_4_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_12_Im = io_in_4_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_13_Re = io_in_13_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_13_Im = io_in_13_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_14_Re = io_in_22_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_14_Im = io_in_22_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_15_Re = io_in_7_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_15_Im = io_in_7_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_16_Re = io_in_16_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_16_Im = io_in_16_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_17_Re = io_in_25_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_17_Im = io_in_25_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_18_Re = io_in_2_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_18_Im = io_in_2_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_19_Re = io_in_11_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_19_Im = io_in_11_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_20_Re = io_in_20_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_20_Im = io_in_20_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_21_Re = io_in_5_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_21_Im = io_in_5_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_22_Re = io_in_14_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_22_Im = io_in_14_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_23_Re = io_in_23_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_23_Im = io_in_23_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_24_Re = io_in_8_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_24_Im = io_in_8_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_25_Re = io_in_17_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_25_Im = io_in_17_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_26_Re = io_in_26_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_26_Im = io_in_26_Im; // @[FFTDesigns.scala 554:17]
endmodule
module PermutationsBasic_1(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_1_Re = io_in_3_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_1_Im = io_in_3_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_2_Re = io_in_6_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_2_Im = io_in_6_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_3_Re = io_in_9_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_3_Im = io_in_9_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_4_Re = io_in_12_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_4_Im = io_in_12_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_5_Re = io_in_15_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_5_Im = io_in_15_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_6_Re = io_in_18_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_6_Im = io_in_18_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_7_Re = io_in_21_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_7_Im = io_in_21_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_8_Re = io_in_24_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_8_Im = io_in_24_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_9_Re = io_in_1_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_9_Im = io_in_1_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_10_Re = io_in_4_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_10_Im = io_in_4_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_11_Re = io_in_7_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_11_Im = io_in_7_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_12_Re = io_in_10_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_12_Im = io_in_10_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_13_Re = io_in_13_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_13_Im = io_in_13_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_14_Re = io_in_16_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_14_Im = io_in_16_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_15_Re = io_in_19_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_15_Im = io_in_19_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_16_Re = io_in_22_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_16_Im = io_in_22_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_17_Re = io_in_25_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_17_Im = io_in_25_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_18_Re = io_in_2_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_18_Im = io_in_2_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_19_Re = io_in_5_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_19_Im = io_in_5_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_20_Re = io_in_8_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_20_Im = io_in_8_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_21_Re = io_in_11_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_21_Im = io_in_11_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_22_Re = io_in_14_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_22_Im = io_in_14_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_23_Re = io_in_17_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_23_Im = io_in_17_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_24_Re = io_in_20_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_24_Im = io_in_20_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_25_Re = io_in_23_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_25_Im = io_in_23_Im; // @[FFTDesigns.scala 554:17]
  assign io_out_26_Re = io_in_26_Re; // @[FFTDesigns.scala 554:17]
  assign io_out_26_Im = io_in_26_Im; // @[FFTDesigns.scala 554:17]
endmodule
module FPComplexMult(
  input         clock,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 45:24]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 45:24]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 45:24]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 45:24]
  wire  FP_adder_clock; // @[FPComplex.scala 46:24]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 46:24]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 46:24]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 46:24]
  wire  FP_multiplier_clock; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 48:26]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 48:26]
  wire  FP_multiplier_2_clock; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_2_io_in_a; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_2_io_in_b; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_2_io_out_s; // @[FPComplex.scala 48:26]
  wire  FP_multiplier_3_clock; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_3_io_in_a; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_3_io_in_b; // @[FPComplex.scala 48:26]
  wire [31:0] FP_multiplier_3_io_out_s; // @[FPComplex.scala 48:26]
  FP_subber FP_subber ( // @[FPComplex.scala 45:24]
    .clock(FP_subber_clock),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 46:24]
    .clock(FP_adder_clock),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 48:26]
    .clock(FP_multiplier_clock),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 48:26]
    .clock(FP_multiplier_1_clock),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  FP_multiplier FP_multiplier_2 ( // @[FPComplex.scala 48:26]
    .clock(FP_multiplier_2_clock),
    .io_in_a(FP_multiplier_2_io_in_a),
    .io_in_b(FP_multiplier_2_io_in_b),
    .io_out_s(FP_multiplier_2_io_out_s)
  );
  FP_multiplier FP_multiplier_3 ( // @[FPComplex.scala 48:26]
    .clock(FP_multiplier_3_clock),
    .io_in_a(FP_multiplier_3_io_in_a),
    .io_in_b(FP_multiplier_3_io_in_b),
    .io_out_s(FP_multiplier_3_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 63:17]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 64:17]
  assign FP_subber_clock = clock;
  assign FP_subber_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 59:17]
  assign FP_subber_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 60:17]
  assign FP_adder_clock = clock;
  assign FP_adder_io_in_a = FP_multiplier_2_io_out_s; // @[FPComplex.scala 61:17]
  assign FP_adder_io_in_b = FP_multiplier_3_io_out_s; // @[FPComplex.scala 62:17]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 51:28]
  assign FP_multiplier_io_in_b = io_in_b_Re; // @[FPComplex.scala 52:28]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 53:28]
  assign FP_multiplier_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 54:28]
  assign FP_multiplier_2_clock = clock;
  assign FP_multiplier_2_io_in_a = io_in_a_Re; // @[FPComplex.scala 55:28]
  assign FP_multiplier_2_io_in_b = io_in_b_Im; // @[FPComplex.scala 56:28]
  assign FP_multiplier_3_clock = clock;
  assign FP_multiplier_3_io_in_a = io_in_a_Im; // @[FPComplex.scala 57:28]
  assign FP_multiplier_3_io_in_b = io_in_b_Re; // @[FPComplex.scala 58:28]
endmodule
module TwiddleFactors(
  input         clock,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_12_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_13_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_14_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_15_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_16_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_17_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_18_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_19_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_20_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_21_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_22_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_23_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_24_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_25_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_26_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  reg [31:0] cnt; // @[FFTDesigns.scala 527:18]
  reg [31:0] cnt2; // @[FFTDesigns.scala 528:19]
  wire [31:0] _cnt_T_1 = cnt + 32'h1; // @[FFTDesigns.scala 534:20]
  wire [31:0] _cnt2_T_1 = cnt2 + 32'h1; // @[FFTDesigns.scala 538:20]
  wire [36:0] _T_2 = cnt * 5'h1b; // @[FFTDesigns.scala 541:58]
  wire [37:0] _T_3 = {{1'd0}, _T_2}; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_13 = 5'ha == _T_3[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_14 = 5'hb == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_13; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_15 = 5'hc == _T_3[4:0] ? 32'h3f800000 : _GEN_14; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_16 = 5'hd == _T_3[4:0] ? 32'h3f441b7c : _GEN_15; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_17 = 5'he == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_16; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_18 = 5'hf == _T_3[4:0] ? 32'h3f800000 : _GEN_17; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_19 = 5'h10 == _T_3[4:0] ? 32'h3f441b7c : _GEN_18; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_20 = 5'h11 == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_19; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_21 = 5'h12 == _T_3[4:0] ? 32'h3f800000 : _GEN_20; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_22 = 5'h13 == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_21; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_23 = 5'h14 == _T_3[4:0] ? 32'hbf708fb2 : _GEN_22; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_24 = 5'h15 == _T_3[4:0] ? 32'h3f800000 : _GEN_23; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_25 = 5'h16 == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_24; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_26 = 5'h17 == _T_3[4:0] ? 32'hbf708fb2 : _GEN_25; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_27 = 5'h18 == _T_3[4:0] ? 32'h3f800000 : _GEN_26; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_28 = 5'h19 == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_27; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_40 = 5'ha == _T_3[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_41 = 5'hb == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_40; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_42 = 5'hc == _T_3[4:0] ? 32'h80800000 : _GEN_41; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_43 = 5'hd == _T_3[4:0] ? 32'hbf248dba : _GEN_42; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_44 = 5'he == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_43; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_45 = 5'hf == _T_3[4:0] ? 32'h80800000 : _GEN_44; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_46 = 5'h10 == _T_3[4:0] ? 32'hbf248dba : _GEN_45; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_47 = 5'h11 == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_46; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_48 = 5'h12 == _T_3[4:0] ? 32'h80800000 : _GEN_47; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_49 = 5'h13 == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_48; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_50 = 5'h14 == _T_3[4:0] ? 32'hbeaf1d40 : _GEN_49; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_51 = 5'h15 == _T_3[4:0] ? 32'h80800000 : _GEN_50; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_52 = 5'h16 == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_51; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_53 = 5'h17 == _T_3[4:0] ? 32'hbeaf1d40 : _GEN_52; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_54 = 5'h18 == _T_3[4:0] ? 32'h80800000 : _GEN_53; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_55 = 5'h19 == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_54; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_58 = 5'h1 == _T_3[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_59 = 5'h2 == _T_3[4:0] ? io_in_2_Im : _GEN_58; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_60 = 5'h3 == _T_3[4:0] ? io_in_3_Im : _GEN_59; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_61 = 5'h4 == _T_3[4:0] ? io_in_4_Im : _GEN_60; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_62 = 5'h5 == _T_3[4:0] ? io_in_5_Im : _GEN_61; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_63 = 5'h6 == _T_3[4:0] ? io_in_6_Im : _GEN_62; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_64 = 5'h7 == _T_3[4:0] ? io_in_7_Im : _GEN_63; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_65 = 5'h8 == _T_3[4:0] ? io_in_8_Im : _GEN_64; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_66 = 5'h9 == _T_3[4:0] ? io_in_9_Im : _GEN_65; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_67 = 5'ha == _T_3[4:0] ? io_in_10_Im : _GEN_66; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_68 = 5'hb == _T_3[4:0] ? io_in_11_Im : _GEN_67; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_69 = 5'hc == _T_3[4:0] ? io_in_12_Im : _GEN_68; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_70 = 5'hd == _T_3[4:0] ? io_in_13_Im : _GEN_69; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_71 = 5'he == _T_3[4:0] ? io_in_14_Im : _GEN_70; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_72 = 5'hf == _T_3[4:0] ? io_in_15_Im : _GEN_71; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_73 = 5'h10 == _T_3[4:0] ? io_in_16_Im : _GEN_72; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_74 = 5'h11 == _T_3[4:0] ? io_in_17_Im : _GEN_73; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_75 = 5'h12 == _T_3[4:0] ? io_in_18_Im : _GEN_74; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_76 = 5'h13 == _T_3[4:0] ? io_in_19_Im : _GEN_75; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_77 = 5'h14 == _T_3[4:0] ? io_in_20_Im : _GEN_76; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_78 = 5'h15 == _T_3[4:0] ? io_in_21_Im : _GEN_77; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_79 = 5'h16 == _T_3[4:0] ? io_in_22_Im : _GEN_78; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_80 = 5'h17 == _T_3[4:0] ? io_in_23_Im : _GEN_79; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_81 = 5'h18 == _T_3[4:0] ? io_in_24_Im : _GEN_80; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_82 = 5'h19 == _T_3[4:0] ? io_in_25_Im : _GEN_81; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_85 = 5'h1 == _T_3[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_86 = 5'h2 == _T_3[4:0] ? io_in_2_Re : _GEN_85; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_87 = 5'h3 == _T_3[4:0] ? io_in_3_Re : _GEN_86; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_88 = 5'h4 == _T_3[4:0] ? io_in_4_Re : _GEN_87; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_89 = 5'h5 == _T_3[4:0] ? io_in_5_Re : _GEN_88; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_90 = 5'h6 == _T_3[4:0] ? io_in_6_Re : _GEN_89; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_91 = 5'h7 == _T_3[4:0] ? io_in_7_Re : _GEN_90; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_92 = 5'h8 == _T_3[4:0] ? io_in_8_Re : _GEN_91; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_93 = 5'h9 == _T_3[4:0] ? io_in_9_Re : _GEN_92; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_94 = 5'ha == _T_3[4:0] ? io_in_10_Re : _GEN_93; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_95 = 5'hb == _T_3[4:0] ? io_in_11_Re : _GEN_94; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_96 = 5'hc == _T_3[4:0] ? io_in_12_Re : _GEN_95; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_97 = 5'hd == _T_3[4:0] ? io_in_13_Re : _GEN_96; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_98 = 5'he == _T_3[4:0] ? io_in_14_Re : _GEN_97; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_99 = 5'hf == _T_3[4:0] ? io_in_15_Re : _GEN_98; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_100 = 5'h10 == _T_3[4:0] ? io_in_16_Re : _GEN_99; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_101 = 5'h11 == _T_3[4:0] ? io_in_17_Re : _GEN_100; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_102 = 5'h12 == _T_3[4:0] ? io_in_18_Re : _GEN_101; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_103 = 5'h13 == _T_3[4:0] ? io_in_19_Re : _GEN_102; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_104 = 5'h14 == _T_3[4:0] ? io_in_20_Re : _GEN_103; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_105 = 5'h15 == _T_3[4:0] ? io_in_21_Re : _GEN_104; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_106 = 5'h16 == _T_3[4:0] ? io_in_22_Re : _GEN_105; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_107 = 5'h17 == _T_3[4:0] ? io_in_23_Re : _GEN_106; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_108 = 5'h18 == _T_3[4:0] ? io_in_24_Re : _GEN_107; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_109 = 5'h19 == _T_3[4:0] ? io_in_25_Re : _GEN_108; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_16 = _T_2 + 37'h1; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_121 = 5'ha == _T_16[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_122 = 5'hb == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_121; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_123 = 5'hc == _T_16[4:0] ? 32'h3f800000 : _GEN_122; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_124 = 5'hd == _T_16[4:0] ? 32'h3f441b7c : _GEN_123; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_125 = 5'he == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_124; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_126 = 5'hf == _T_16[4:0] ? 32'h3f800000 : _GEN_125; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_127 = 5'h10 == _T_16[4:0] ? 32'h3f441b7c : _GEN_126; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_128 = 5'h11 == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_127; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_129 = 5'h12 == _T_16[4:0] ? 32'h3f800000 : _GEN_128; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_130 = 5'h13 == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_129; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_131 = 5'h14 == _T_16[4:0] ? 32'hbf708fb2 : _GEN_130; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_132 = 5'h15 == _T_16[4:0] ? 32'h3f800000 : _GEN_131; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_133 = 5'h16 == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_132; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_134 = 5'h17 == _T_16[4:0] ? 32'hbf708fb2 : _GEN_133; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_135 = 5'h18 == _T_16[4:0] ? 32'h3f800000 : _GEN_134; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_136 = 5'h19 == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_135; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_148 = 5'ha == _T_16[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_149 = 5'hb == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_148; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_150 = 5'hc == _T_16[4:0] ? 32'h80800000 : _GEN_149; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_151 = 5'hd == _T_16[4:0] ? 32'hbf248dba : _GEN_150; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_152 = 5'he == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_151; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_153 = 5'hf == _T_16[4:0] ? 32'h80800000 : _GEN_152; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_154 = 5'h10 == _T_16[4:0] ? 32'hbf248dba : _GEN_153; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_155 = 5'h11 == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_154; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_156 = 5'h12 == _T_16[4:0] ? 32'h80800000 : _GEN_155; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_157 = 5'h13 == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_156; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_158 = 5'h14 == _T_16[4:0] ? 32'hbeaf1d40 : _GEN_157; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_159 = 5'h15 == _T_16[4:0] ? 32'h80800000 : _GEN_158; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_160 = 5'h16 == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_159; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_161 = 5'h17 == _T_16[4:0] ? 32'hbeaf1d40 : _GEN_160; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_162 = 5'h18 == _T_16[4:0] ? 32'h80800000 : _GEN_161; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_163 = 5'h19 == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_162; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_166 = 5'h1 == _T_16[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_167 = 5'h2 == _T_16[4:0] ? io_in_2_Im : _GEN_166; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_168 = 5'h3 == _T_16[4:0] ? io_in_3_Im : _GEN_167; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_169 = 5'h4 == _T_16[4:0] ? io_in_4_Im : _GEN_168; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_170 = 5'h5 == _T_16[4:0] ? io_in_5_Im : _GEN_169; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_171 = 5'h6 == _T_16[4:0] ? io_in_6_Im : _GEN_170; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_172 = 5'h7 == _T_16[4:0] ? io_in_7_Im : _GEN_171; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_173 = 5'h8 == _T_16[4:0] ? io_in_8_Im : _GEN_172; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_174 = 5'h9 == _T_16[4:0] ? io_in_9_Im : _GEN_173; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_175 = 5'ha == _T_16[4:0] ? io_in_10_Im : _GEN_174; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_176 = 5'hb == _T_16[4:0] ? io_in_11_Im : _GEN_175; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_177 = 5'hc == _T_16[4:0] ? io_in_12_Im : _GEN_176; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_178 = 5'hd == _T_16[4:0] ? io_in_13_Im : _GEN_177; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_179 = 5'he == _T_16[4:0] ? io_in_14_Im : _GEN_178; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_180 = 5'hf == _T_16[4:0] ? io_in_15_Im : _GEN_179; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_181 = 5'h10 == _T_16[4:0] ? io_in_16_Im : _GEN_180; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_182 = 5'h11 == _T_16[4:0] ? io_in_17_Im : _GEN_181; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_183 = 5'h12 == _T_16[4:0] ? io_in_18_Im : _GEN_182; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_184 = 5'h13 == _T_16[4:0] ? io_in_19_Im : _GEN_183; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_185 = 5'h14 == _T_16[4:0] ? io_in_20_Im : _GEN_184; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_186 = 5'h15 == _T_16[4:0] ? io_in_21_Im : _GEN_185; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_187 = 5'h16 == _T_16[4:0] ? io_in_22_Im : _GEN_186; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_188 = 5'h17 == _T_16[4:0] ? io_in_23_Im : _GEN_187; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_189 = 5'h18 == _T_16[4:0] ? io_in_24_Im : _GEN_188; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_190 = 5'h19 == _T_16[4:0] ? io_in_25_Im : _GEN_189; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_193 = 5'h1 == _T_16[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_194 = 5'h2 == _T_16[4:0] ? io_in_2_Re : _GEN_193; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_195 = 5'h3 == _T_16[4:0] ? io_in_3_Re : _GEN_194; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_196 = 5'h4 == _T_16[4:0] ? io_in_4_Re : _GEN_195; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_197 = 5'h5 == _T_16[4:0] ? io_in_5_Re : _GEN_196; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_198 = 5'h6 == _T_16[4:0] ? io_in_6_Re : _GEN_197; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_199 = 5'h7 == _T_16[4:0] ? io_in_7_Re : _GEN_198; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_200 = 5'h8 == _T_16[4:0] ? io_in_8_Re : _GEN_199; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_201 = 5'h9 == _T_16[4:0] ? io_in_9_Re : _GEN_200; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_202 = 5'ha == _T_16[4:0] ? io_in_10_Re : _GEN_201; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_203 = 5'hb == _T_16[4:0] ? io_in_11_Re : _GEN_202; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_204 = 5'hc == _T_16[4:0] ? io_in_12_Re : _GEN_203; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_205 = 5'hd == _T_16[4:0] ? io_in_13_Re : _GEN_204; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_206 = 5'he == _T_16[4:0] ? io_in_14_Re : _GEN_205; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_207 = 5'hf == _T_16[4:0] ? io_in_15_Re : _GEN_206; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_208 = 5'h10 == _T_16[4:0] ? io_in_16_Re : _GEN_207; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_209 = 5'h11 == _T_16[4:0] ? io_in_17_Re : _GEN_208; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_210 = 5'h12 == _T_16[4:0] ? io_in_18_Re : _GEN_209; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_211 = 5'h13 == _T_16[4:0] ? io_in_19_Re : _GEN_210; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_212 = 5'h14 == _T_16[4:0] ? io_in_20_Re : _GEN_211; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_213 = 5'h15 == _T_16[4:0] ? io_in_21_Re : _GEN_212; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_214 = 5'h16 == _T_16[4:0] ? io_in_22_Re : _GEN_213; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_215 = 5'h17 == _T_16[4:0] ? io_in_23_Re : _GEN_214; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_216 = 5'h18 == _T_16[4:0] ? io_in_24_Re : _GEN_215; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_217 = 5'h19 == _T_16[4:0] ? io_in_25_Re : _GEN_216; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_28 = _T_2 + 37'h2; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_229 = 5'ha == _T_28[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_230 = 5'hb == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_229; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_231 = 5'hc == _T_28[4:0] ? 32'h3f800000 : _GEN_230; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_232 = 5'hd == _T_28[4:0] ? 32'h3f441b7c : _GEN_231; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_233 = 5'he == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_232; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_234 = 5'hf == _T_28[4:0] ? 32'h3f800000 : _GEN_233; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_235 = 5'h10 == _T_28[4:0] ? 32'h3f441b7c : _GEN_234; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_236 = 5'h11 == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_235; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_237 = 5'h12 == _T_28[4:0] ? 32'h3f800000 : _GEN_236; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_238 = 5'h13 == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_237; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_239 = 5'h14 == _T_28[4:0] ? 32'hbf708fb2 : _GEN_238; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_240 = 5'h15 == _T_28[4:0] ? 32'h3f800000 : _GEN_239; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_241 = 5'h16 == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_240; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_242 = 5'h17 == _T_28[4:0] ? 32'hbf708fb2 : _GEN_241; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_243 = 5'h18 == _T_28[4:0] ? 32'h3f800000 : _GEN_242; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_244 = 5'h19 == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_243; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_256 = 5'ha == _T_28[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_257 = 5'hb == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_256; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_258 = 5'hc == _T_28[4:0] ? 32'h80800000 : _GEN_257; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_259 = 5'hd == _T_28[4:0] ? 32'hbf248dba : _GEN_258; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_260 = 5'he == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_259; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_261 = 5'hf == _T_28[4:0] ? 32'h80800000 : _GEN_260; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_262 = 5'h10 == _T_28[4:0] ? 32'hbf248dba : _GEN_261; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_263 = 5'h11 == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_262; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_264 = 5'h12 == _T_28[4:0] ? 32'h80800000 : _GEN_263; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_265 = 5'h13 == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_264; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_266 = 5'h14 == _T_28[4:0] ? 32'hbeaf1d40 : _GEN_265; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_267 = 5'h15 == _T_28[4:0] ? 32'h80800000 : _GEN_266; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_268 = 5'h16 == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_267; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_269 = 5'h17 == _T_28[4:0] ? 32'hbeaf1d40 : _GEN_268; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_270 = 5'h18 == _T_28[4:0] ? 32'h80800000 : _GEN_269; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_271 = 5'h19 == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_270; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_274 = 5'h1 == _T_28[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_275 = 5'h2 == _T_28[4:0] ? io_in_2_Im : _GEN_274; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_276 = 5'h3 == _T_28[4:0] ? io_in_3_Im : _GEN_275; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_277 = 5'h4 == _T_28[4:0] ? io_in_4_Im : _GEN_276; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_278 = 5'h5 == _T_28[4:0] ? io_in_5_Im : _GEN_277; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_279 = 5'h6 == _T_28[4:0] ? io_in_6_Im : _GEN_278; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_280 = 5'h7 == _T_28[4:0] ? io_in_7_Im : _GEN_279; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_281 = 5'h8 == _T_28[4:0] ? io_in_8_Im : _GEN_280; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_282 = 5'h9 == _T_28[4:0] ? io_in_9_Im : _GEN_281; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_283 = 5'ha == _T_28[4:0] ? io_in_10_Im : _GEN_282; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_284 = 5'hb == _T_28[4:0] ? io_in_11_Im : _GEN_283; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_285 = 5'hc == _T_28[4:0] ? io_in_12_Im : _GEN_284; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_286 = 5'hd == _T_28[4:0] ? io_in_13_Im : _GEN_285; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_287 = 5'he == _T_28[4:0] ? io_in_14_Im : _GEN_286; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_288 = 5'hf == _T_28[4:0] ? io_in_15_Im : _GEN_287; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_289 = 5'h10 == _T_28[4:0] ? io_in_16_Im : _GEN_288; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_290 = 5'h11 == _T_28[4:0] ? io_in_17_Im : _GEN_289; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_291 = 5'h12 == _T_28[4:0] ? io_in_18_Im : _GEN_290; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_292 = 5'h13 == _T_28[4:0] ? io_in_19_Im : _GEN_291; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_293 = 5'h14 == _T_28[4:0] ? io_in_20_Im : _GEN_292; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_294 = 5'h15 == _T_28[4:0] ? io_in_21_Im : _GEN_293; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_295 = 5'h16 == _T_28[4:0] ? io_in_22_Im : _GEN_294; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_296 = 5'h17 == _T_28[4:0] ? io_in_23_Im : _GEN_295; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_297 = 5'h18 == _T_28[4:0] ? io_in_24_Im : _GEN_296; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_298 = 5'h19 == _T_28[4:0] ? io_in_25_Im : _GEN_297; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_301 = 5'h1 == _T_28[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_302 = 5'h2 == _T_28[4:0] ? io_in_2_Re : _GEN_301; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_303 = 5'h3 == _T_28[4:0] ? io_in_3_Re : _GEN_302; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_304 = 5'h4 == _T_28[4:0] ? io_in_4_Re : _GEN_303; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_305 = 5'h5 == _T_28[4:0] ? io_in_5_Re : _GEN_304; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_306 = 5'h6 == _T_28[4:0] ? io_in_6_Re : _GEN_305; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_307 = 5'h7 == _T_28[4:0] ? io_in_7_Re : _GEN_306; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_308 = 5'h8 == _T_28[4:0] ? io_in_8_Re : _GEN_307; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_309 = 5'h9 == _T_28[4:0] ? io_in_9_Re : _GEN_308; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_310 = 5'ha == _T_28[4:0] ? io_in_10_Re : _GEN_309; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_311 = 5'hb == _T_28[4:0] ? io_in_11_Re : _GEN_310; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_312 = 5'hc == _T_28[4:0] ? io_in_12_Re : _GEN_311; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_313 = 5'hd == _T_28[4:0] ? io_in_13_Re : _GEN_312; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_314 = 5'he == _T_28[4:0] ? io_in_14_Re : _GEN_313; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_315 = 5'hf == _T_28[4:0] ? io_in_15_Re : _GEN_314; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_316 = 5'h10 == _T_28[4:0] ? io_in_16_Re : _GEN_315; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_317 = 5'h11 == _T_28[4:0] ? io_in_17_Re : _GEN_316; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_318 = 5'h12 == _T_28[4:0] ? io_in_18_Re : _GEN_317; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_319 = 5'h13 == _T_28[4:0] ? io_in_19_Re : _GEN_318; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_320 = 5'h14 == _T_28[4:0] ? io_in_20_Re : _GEN_319; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_321 = 5'h15 == _T_28[4:0] ? io_in_21_Re : _GEN_320; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_322 = 5'h16 == _T_28[4:0] ? io_in_22_Re : _GEN_321; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_323 = 5'h17 == _T_28[4:0] ? io_in_23_Re : _GEN_322; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_324 = 5'h18 == _T_28[4:0] ? io_in_24_Re : _GEN_323; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_325 = 5'h19 == _T_28[4:0] ? io_in_25_Re : _GEN_324; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_40 = _T_2 + 37'h3; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_337 = 5'ha == _T_40[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_338 = 5'hb == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_337; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_339 = 5'hc == _T_40[4:0] ? 32'h3f800000 : _GEN_338; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_340 = 5'hd == _T_40[4:0] ? 32'h3f441b7c : _GEN_339; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_341 = 5'he == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_340; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_342 = 5'hf == _T_40[4:0] ? 32'h3f800000 : _GEN_341; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_343 = 5'h10 == _T_40[4:0] ? 32'h3f441b7c : _GEN_342; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_344 = 5'h11 == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_343; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_345 = 5'h12 == _T_40[4:0] ? 32'h3f800000 : _GEN_344; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_346 = 5'h13 == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_345; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_347 = 5'h14 == _T_40[4:0] ? 32'hbf708fb2 : _GEN_346; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_348 = 5'h15 == _T_40[4:0] ? 32'h3f800000 : _GEN_347; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_349 = 5'h16 == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_348; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_350 = 5'h17 == _T_40[4:0] ? 32'hbf708fb2 : _GEN_349; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_351 = 5'h18 == _T_40[4:0] ? 32'h3f800000 : _GEN_350; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_352 = 5'h19 == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_351; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_364 = 5'ha == _T_40[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_365 = 5'hb == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_364; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_366 = 5'hc == _T_40[4:0] ? 32'h80800000 : _GEN_365; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_367 = 5'hd == _T_40[4:0] ? 32'hbf248dba : _GEN_366; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_368 = 5'he == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_367; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_369 = 5'hf == _T_40[4:0] ? 32'h80800000 : _GEN_368; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_370 = 5'h10 == _T_40[4:0] ? 32'hbf248dba : _GEN_369; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_371 = 5'h11 == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_370; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_372 = 5'h12 == _T_40[4:0] ? 32'h80800000 : _GEN_371; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_373 = 5'h13 == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_372; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_374 = 5'h14 == _T_40[4:0] ? 32'hbeaf1d40 : _GEN_373; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_375 = 5'h15 == _T_40[4:0] ? 32'h80800000 : _GEN_374; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_376 = 5'h16 == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_375; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_377 = 5'h17 == _T_40[4:0] ? 32'hbeaf1d40 : _GEN_376; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_378 = 5'h18 == _T_40[4:0] ? 32'h80800000 : _GEN_377; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_379 = 5'h19 == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_378; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_382 = 5'h1 == _T_40[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_383 = 5'h2 == _T_40[4:0] ? io_in_2_Im : _GEN_382; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_384 = 5'h3 == _T_40[4:0] ? io_in_3_Im : _GEN_383; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_385 = 5'h4 == _T_40[4:0] ? io_in_4_Im : _GEN_384; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_386 = 5'h5 == _T_40[4:0] ? io_in_5_Im : _GEN_385; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_387 = 5'h6 == _T_40[4:0] ? io_in_6_Im : _GEN_386; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_388 = 5'h7 == _T_40[4:0] ? io_in_7_Im : _GEN_387; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_389 = 5'h8 == _T_40[4:0] ? io_in_8_Im : _GEN_388; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_390 = 5'h9 == _T_40[4:0] ? io_in_9_Im : _GEN_389; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_391 = 5'ha == _T_40[4:0] ? io_in_10_Im : _GEN_390; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_392 = 5'hb == _T_40[4:0] ? io_in_11_Im : _GEN_391; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_393 = 5'hc == _T_40[4:0] ? io_in_12_Im : _GEN_392; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_394 = 5'hd == _T_40[4:0] ? io_in_13_Im : _GEN_393; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_395 = 5'he == _T_40[4:0] ? io_in_14_Im : _GEN_394; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_396 = 5'hf == _T_40[4:0] ? io_in_15_Im : _GEN_395; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_397 = 5'h10 == _T_40[4:0] ? io_in_16_Im : _GEN_396; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_398 = 5'h11 == _T_40[4:0] ? io_in_17_Im : _GEN_397; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_399 = 5'h12 == _T_40[4:0] ? io_in_18_Im : _GEN_398; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_400 = 5'h13 == _T_40[4:0] ? io_in_19_Im : _GEN_399; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_401 = 5'h14 == _T_40[4:0] ? io_in_20_Im : _GEN_400; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_402 = 5'h15 == _T_40[4:0] ? io_in_21_Im : _GEN_401; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_403 = 5'h16 == _T_40[4:0] ? io_in_22_Im : _GEN_402; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_404 = 5'h17 == _T_40[4:0] ? io_in_23_Im : _GEN_403; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_405 = 5'h18 == _T_40[4:0] ? io_in_24_Im : _GEN_404; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_406 = 5'h19 == _T_40[4:0] ? io_in_25_Im : _GEN_405; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_409 = 5'h1 == _T_40[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_410 = 5'h2 == _T_40[4:0] ? io_in_2_Re : _GEN_409; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_411 = 5'h3 == _T_40[4:0] ? io_in_3_Re : _GEN_410; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_412 = 5'h4 == _T_40[4:0] ? io_in_4_Re : _GEN_411; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_413 = 5'h5 == _T_40[4:0] ? io_in_5_Re : _GEN_412; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_414 = 5'h6 == _T_40[4:0] ? io_in_6_Re : _GEN_413; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_415 = 5'h7 == _T_40[4:0] ? io_in_7_Re : _GEN_414; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_416 = 5'h8 == _T_40[4:0] ? io_in_8_Re : _GEN_415; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_417 = 5'h9 == _T_40[4:0] ? io_in_9_Re : _GEN_416; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_418 = 5'ha == _T_40[4:0] ? io_in_10_Re : _GEN_417; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_419 = 5'hb == _T_40[4:0] ? io_in_11_Re : _GEN_418; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_420 = 5'hc == _T_40[4:0] ? io_in_12_Re : _GEN_419; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_421 = 5'hd == _T_40[4:0] ? io_in_13_Re : _GEN_420; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_422 = 5'he == _T_40[4:0] ? io_in_14_Re : _GEN_421; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_423 = 5'hf == _T_40[4:0] ? io_in_15_Re : _GEN_422; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_424 = 5'h10 == _T_40[4:0] ? io_in_16_Re : _GEN_423; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_425 = 5'h11 == _T_40[4:0] ? io_in_17_Re : _GEN_424; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_426 = 5'h12 == _T_40[4:0] ? io_in_18_Re : _GEN_425; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_427 = 5'h13 == _T_40[4:0] ? io_in_19_Re : _GEN_426; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_428 = 5'h14 == _T_40[4:0] ? io_in_20_Re : _GEN_427; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_429 = 5'h15 == _T_40[4:0] ? io_in_21_Re : _GEN_428; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_430 = 5'h16 == _T_40[4:0] ? io_in_22_Re : _GEN_429; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_431 = 5'h17 == _T_40[4:0] ? io_in_23_Re : _GEN_430; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_432 = 5'h18 == _T_40[4:0] ? io_in_24_Re : _GEN_431; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_433 = 5'h19 == _T_40[4:0] ? io_in_25_Re : _GEN_432; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_52 = _T_2 + 37'h4; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_445 = 5'ha == _T_52[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_446 = 5'hb == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_445; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_447 = 5'hc == _T_52[4:0] ? 32'h3f800000 : _GEN_446; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_448 = 5'hd == _T_52[4:0] ? 32'h3f441b7c : _GEN_447; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_449 = 5'he == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_448; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_450 = 5'hf == _T_52[4:0] ? 32'h3f800000 : _GEN_449; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_451 = 5'h10 == _T_52[4:0] ? 32'h3f441b7c : _GEN_450; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_452 = 5'h11 == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_451; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_453 = 5'h12 == _T_52[4:0] ? 32'h3f800000 : _GEN_452; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_454 = 5'h13 == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_453; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_455 = 5'h14 == _T_52[4:0] ? 32'hbf708fb2 : _GEN_454; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_456 = 5'h15 == _T_52[4:0] ? 32'h3f800000 : _GEN_455; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_457 = 5'h16 == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_456; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_458 = 5'h17 == _T_52[4:0] ? 32'hbf708fb2 : _GEN_457; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_459 = 5'h18 == _T_52[4:0] ? 32'h3f800000 : _GEN_458; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_460 = 5'h19 == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_459; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_472 = 5'ha == _T_52[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_473 = 5'hb == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_472; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_474 = 5'hc == _T_52[4:0] ? 32'h80800000 : _GEN_473; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_475 = 5'hd == _T_52[4:0] ? 32'hbf248dba : _GEN_474; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_476 = 5'he == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_475; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_477 = 5'hf == _T_52[4:0] ? 32'h80800000 : _GEN_476; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_478 = 5'h10 == _T_52[4:0] ? 32'hbf248dba : _GEN_477; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_479 = 5'h11 == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_478; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_480 = 5'h12 == _T_52[4:0] ? 32'h80800000 : _GEN_479; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_481 = 5'h13 == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_480; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_482 = 5'h14 == _T_52[4:0] ? 32'hbeaf1d40 : _GEN_481; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_483 = 5'h15 == _T_52[4:0] ? 32'h80800000 : _GEN_482; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_484 = 5'h16 == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_483; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_485 = 5'h17 == _T_52[4:0] ? 32'hbeaf1d40 : _GEN_484; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_486 = 5'h18 == _T_52[4:0] ? 32'h80800000 : _GEN_485; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_487 = 5'h19 == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_486; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_490 = 5'h1 == _T_52[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_491 = 5'h2 == _T_52[4:0] ? io_in_2_Im : _GEN_490; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_492 = 5'h3 == _T_52[4:0] ? io_in_3_Im : _GEN_491; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_493 = 5'h4 == _T_52[4:0] ? io_in_4_Im : _GEN_492; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_494 = 5'h5 == _T_52[4:0] ? io_in_5_Im : _GEN_493; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_495 = 5'h6 == _T_52[4:0] ? io_in_6_Im : _GEN_494; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_496 = 5'h7 == _T_52[4:0] ? io_in_7_Im : _GEN_495; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_497 = 5'h8 == _T_52[4:0] ? io_in_8_Im : _GEN_496; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_498 = 5'h9 == _T_52[4:0] ? io_in_9_Im : _GEN_497; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_499 = 5'ha == _T_52[4:0] ? io_in_10_Im : _GEN_498; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_500 = 5'hb == _T_52[4:0] ? io_in_11_Im : _GEN_499; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_501 = 5'hc == _T_52[4:0] ? io_in_12_Im : _GEN_500; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_502 = 5'hd == _T_52[4:0] ? io_in_13_Im : _GEN_501; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_503 = 5'he == _T_52[4:0] ? io_in_14_Im : _GEN_502; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_504 = 5'hf == _T_52[4:0] ? io_in_15_Im : _GEN_503; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_505 = 5'h10 == _T_52[4:0] ? io_in_16_Im : _GEN_504; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_506 = 5'h11 == _T_52[4:0] ? io_in_17_Im : _GEN_505; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_507 = 5'h12 == _T_52[4:0] ? io_in_18_Im : _GEN_506; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_508 = 5'h13 == _T_52[4:0] ? io_in_19_Im : _GEN_507; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_509 = 5'h14 == _T_52[4:0] ? io_in_20_Im : _GEN_508; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_510 = 5'h15 == _T_52[4:0] ? io_in_21_Im : _GEN_509; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_511 = 5'h16 == _T_52[4:0] ? io_in_22_Im : _GEN_510; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_512 = 5'h17 == _T_52[4:0] ? io_in_23_Im : _GEN_511; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_513 = 5'h18 == _T_52[4:0] ? io_in_24_Im : _GEN_512; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_514 = 5'h19 == _T_52[4:0] ? io_in_25_Im : _GEN_513; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_517 = 5'h1 == _T_52[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_518 = 5'h2 == _T_52[4:0] ? io_in_2_Re : _GEN_517; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_519 = 5'h3 == _T_52[4:0] ? io_in_3_Re : _GEN_518; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_520 = 5'h4 == _T_52[4:0] ? io_in_4_Re : _GEN_519; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_521 = 5'h5 == _T_52[4:0] ? io_in_5_Re : _GEN_520; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_522 = 5'h6 == _T_52[4:0] ? io_in_6_Re : _GEN_521; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_523 = 5'h7 == _T_52[4:0] ? io_in_7_Re : _GEN_522; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_524 = 5'h8 == _T_52[4:0] ? io_in_8_Re : _GEN_523; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_525 = 5'h9 == _T_52[4:0] ? io_in_9_Re : _GEN_524; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_526 = 5'ha == _T_52[4:0] ? io_in_10_Re : _GEN_525; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_527 = 5'hb == _T_52[4:0] ? io_in_11_Re : _GEN_526; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_528 = 5'hc == _T_52[4:0] ? io_in_12_Re : _GEN_527; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_529 = 5'hd == _T_52[4:0] ? io_in_13_Re : _GEN_528; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_530 = 5'he == _T_52[4:0] ? io_in_14_Re : _GEN_529; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_531 = 5'hf == _T_52[4:0] ? io_in_15_Re : _GEN_530; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_532 = 5'h10 == _T_52[4:0] ? io_in_16_Re : _GEN_531; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_533 = 5'h11 == _T_52[4:0] ? io_in_17_Re : _GEN_532; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_534 = 5'h12 == _T_52[4:0] ? io_in_18_Re : _GEN_533; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_535 = 5'h13 == _T_52[4:0] ? io_in_19_Re : _GEN_534; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_536 = 5'h14 == _T_52[4:0] ? io_in_20_Re : _GEN_535; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_537 = 5'h15 == _T_52[4:0] ? io_in_21_Re : _GEN_536; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_538 = 5'h16 == _T_52[4:0] ? io_in_22_Re : _GEN_537; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_539 = 5'h17 == _T_52[4:0] ? io_in_23_Re : _GEN_538; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_540 = 5'h18 == _T_52[4:0] ? io_in_24_Re : _GEN_539; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_541 = 5'h19 == _T_52[4:0] ? io_in_25_Re : _GEN_540; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_64 = _T_2 + 37'h5; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_553 = 5'ha == _T_64[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_554 = 5'hb == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_553; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_555 = 5'hc == _T_64[4:0] ? 32'h3f800000 : _GEN_554; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_556 = 5'hd == _T_64[4:0] ? 32'h3f441b7c : _GEN_555; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_557 = 5'he == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_556; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_558 = 5'hf == _T_64[4:0] ? 32'h3f800000 : _GEN_557; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_559 = 5'h10 == _T_64[4:0] ? 32'h3f441b7c : _GEN_558; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_560 = 5'h11 == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_559; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_561 = 5'h12 == _T_64[4:0] ? 32'h3f800000 : _GEN_560; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_562 = 5'h13 == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_561; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_563 = 5'h14 == _T_64[4:0] ? 32'hbf708fb2 : _GEN_562; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_564 = 5'h15 == _T_64[4:0] ? 32'h3f800000 : _GEN_563; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_565 = 5'h16 == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_564; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_566 = 5'h17 == _T_64[4:0] ? 32'hbf708fb2 : _GEN_565; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_567 = 5'h18 == _T_64[4:0] ? 32'h3f800000 : _GEN_566; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_568 = 5'h19 == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_567; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_580 = 5'ha == _T_64[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_581 = 5'hb == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_580; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_582 = 5'hc == _T_64[4:0] ? 32'h80800000 : _GEN_581; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_583 = 5'hd == _T_64[4:0] ? 32'hbf248dba : _GEN_582; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_584 = 5'he == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_583; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_585 = 5'hf == _T_64[4:0] ? 32'h80800000 : _GEN_584; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_586 = 5'h10 == _T_64[4:0] ? 32'hbf248dba : _GEN_585; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_587 = 5'h11 == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_586; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_588 = 5'h12 == _T_64[4:0] ? 32'h80800000 : _GEN_587; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_589 = 5'h13 == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_588; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_590 = 5'h14 == _T_64[4:0] ? 32'hbeaf1d40 : _GEN_589; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_591 = 5'h15 == _T_64[4:0] ? 32'h80800000 : _GEN_590; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_592 = 5'h16 == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_591; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_593 = 5'h17 == _T_64[4:0] ? 32'hbeaf1d40 : _GEN_592; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_594 = 5'h18 == _T_64[4:0] ? 32'h80800000 : _GEN_593; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_595 = 5'h19 == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_594; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_598 = 5'h1 == _T_64[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_599 = 5'h2 == _T_64[4:0] ? io_in_2_Im : _GEN_598; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_600 = 5'h3 == _T_64[4:0] ? io_in_3_Im : _GEN_599; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_601 = 5'h4 == _T_64[4:0] ? io_in_4_Im : _GEN_600; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_602 = 5'h5 == _T_64[4:0] ? io_in_5_Im : _GEN_601; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_603 = 5'h6 == _T_64[4:0] ? io_in_6_Im : _GEN_602; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_604 = 5'h7 == _T_64[4:0] ? io_in_7_Im : _GEN_603; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_605 = 5'h8 == _T_64[4:0] ? io_in_8_Im : _GEN_604; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_606 = 5'h9 == _T_64[4:0] ? io_in_9_Im : _GEN_605; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_607 = 5'ha == _T_64[4:0] ? io_in_10_Im : _GEN_606; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_608 = 5'hb == _T_64[4:0] ? io_in_11_Im : _GEN_607; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_609 = 5'hc == _T_64[4:0] ? io_in_12_Im : _GEN_608; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_610 = 5'hd == _T_64[4:0] ? io_in_13_Im : _GEN_609; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_611 = 5'he == _T_64[4:0] ? io_in_14_Im : _GEN_610; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_612 = 5'hf == _T_64[4:0] ? io_in_15_Im : _GEN_611; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_613 = 5'h10 == _T_64[4:0] ? io_in_16_Im : _GEN_612; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_614 = 5'h11 == _T_64[4:0] ? io_in_17_Im : _GEN_613; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_615 = 5'h12 == _T_64[4:0] ? io_in_18_Im : _GEN_614; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_616 = 5'h13 == _T_64[4:0] ? io_in_19_Im : _GEN_615; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_617 = 5'h14 == _T_64[4:0] ? io_in_20_Im : _GEN_616; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_618 = 5'h15 == _T_64[4:0] ? io_in_21_Im : _GEN_617; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_619 = 5'h16 == _T_64[4:0] ? io_in_22_Im : _GEN_618; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_620 = 5'h17 == _T_64[4:0] ? io_in_23_Im : _GEN_619; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_621 = 5'h18 == _T_64[4:0] ? io_in_24_Im : _GEN_620; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_622 = 5'h19 == _T_64[4:0] ? io_in_25_Im : _GEN_621; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_625 = 5'h1 == _T_64[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_626 = 5'h2 == _T_64[4:0] ? io_in_2_Re : _GEN_625; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_627 = 5'h3 == _T_64[4:0] ? io_in_3_Re : _GEN_626; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_628 = 5'h4 == _T_64[4:0] ? io_in_4_Re : _GEN_627; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_629 = 5'h5 == _T_64[4:0] ? io_in_5_Re : _GEN_628; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_630 = 5'h6 == _T_64[4:0] ? io_in_6_Re : _GEN_629; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_631 = 5'h7 == _T_64[4:0] ? io_in_7_Re : _GEN_630; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_632 = 5'h8 == _T_64[4:0] ? io_in_8_Re : _GEN_631; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_633 = 5'h9 == _T_64[4:0] ? io_in_9_Re : _GEN_632; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_634 = 5'ha == _T_64[4:0] ? io_in_10_Re : _GEN_633; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_635 = 5'hb == _T_64[4:0] ? io_in_11_Re : _GEN_634; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_636 = 5'hc == _T_64[4:0] ? io_in_12_Re : _GEN_635; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_637 = 5'hd == _T_64[4:0] ? io_in_13_Re : _GEN_636; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_638 = 5'he == _T_64[4:0] ? io_in_14_Re : _GEN_637; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_639 = 5'hf == _T_64[4:0] ? io_in_15_Re : _GEN_638; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_640 = 5'h10 == _T_64[4:0] ? io_in_16_Re : _GEN_639; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_641 = 5'h11 == _T_64[4:0] ? io_in_17_Re : _GEN_640; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_642 = 5'h12 == _T_64[4:0] ? io_in_18_Re : _GEN_641; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_643 = 5'h13 == _T_64[4:0] ? io_in_19_Re : _GEN_642; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_644 = 5'h14 == _T_64[4:0] ? io_in_20_Re : _GEN_643; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_645 = 5'h15 == _T_64[4:0] ? io_in_21_Re : _GEN_644; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_646 = 5'h16 == _T_64[4:0] ? io_in_22_Re : _GEN_645; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_647 = 5'h17 == _T_64[4:0] ? io_in_23_Re : _GEN_646; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_648 = 5'h18 == _T_64[4:0] ? io_in_24_Re : _GEN_647; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_649 = 5'h19 == _T_64[4:0] ? io_in_25_Re : _GEN_648; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_76 = _T_2 + 37'h6; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_661 = 5'ha == _T_76[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_662 = 5'hb == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_661; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_663 = 5'hc == _T_76[4:0] ? 32'h3f800000 : _GEN_662; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_664 = 5'hd == _T_76[4:0] ? 32'h3f441b7c : _GEN_663; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_665 = 5'he == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_664; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_666 = 5'hf == _T_76[4:0] ? 32'h3f800000 : _GEN_665; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_667 = 5'h10 == _T_76[4:0] ? 32'h3f441b7c : _GEN_666; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_668 = 5'h11 == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_667; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_669 = 5'h12 == _T_76[4:0] ? 32'h3f800000 : _GEN_668; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_670 = 5'h13 == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_669; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_671 = 5'h14 == _T_76[4:0] ? 32'hbf708fb2 : _GEN_670; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_672 = 5'h15 == _T_76[4:0] ? 32'h3f800000 : _GEN_671; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_673 = 5'h16 == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_672; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_674 = 5'h17 == _T_76[4:0] ? 32'hbf708fb2 : _GEN_673; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_675 = 5'h18 == _T_76[4:0] ? 32'h3f800000 : _GEN_674; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_676 = 5'h19 == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_675; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_688 = 5'ha == _T_76[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_689 = 5'hb == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_688; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_690 = 5'hc == _T_76[4:0] ? 32'h80800000 : _GEN_689; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_691 = 5'hd == _T_76[4:0] ? 32'hbf248dba : _GEN_690; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_692 = 5'he == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_691; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_693 = 5'hf == _T_76[4:0] ? 32'h80800000 : _GEN_692; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_694 = 5'h10 == _T_76[4:0] ? 32'hbf248dba : _GEN_693; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_695 = 5'h11 == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_694; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_696 = 5'h12 == _T_76[4:0] ? 32'h80800000 : _GEN_695; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_697 = 5'h13 == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_696; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_698 = 5'h14 == _T_76[4:0] ? 32'hbeaf1d40 : _GEN_697; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_699 = 5'h15 == _T_76[4:0] ? 32'h80800000 : _GEN_698; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_700 = 5'h16 == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_699; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_701 = 5'h17 == _T_76[4:0] ? 32'hbeaf1d40 : _GEN_700; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_702 = 5'h18 == _T_76[4:0] ? 32'h80800000 : _GEN_701; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_703 = 5'h19 == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_702; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_706 = 5'h1 == _T_76[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_707 = 5'h2 == _T_76[4:0] ? io_in_2_Im : _GEN_706; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_708 = 5'h3 == _T_76[4:0] ? io_in_3_Im : _GEN_707; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_709 = 5'h4 == _T_76[4:0] ? io_in_4_Im : _GEN_708; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_710 = 5'h5 == _T_76[4:0] ? io_in_5_Im : _GEN_709; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_711 = 5'h6 == _T_76[4:0] ? io_in_6_Im : _GEN_710; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_712 = 5'h7 == _T_76[4:0] ? io_in_7_Im : _GEN_711; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_713 = 5'h8 == _T_76[4:0] ? io_in_8_Im : _GEN_712; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_714 = 5'h9 == _T_76[4:0] ? io_in_9_Im : _GEN_713; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_715 = 5'ha == _T_76[4:0] ? io_in_10_Im : _GEN_714; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_716 = 5'hb == _T_76[4:0] ? io_in_11_Im : _GEN_715; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_717 = 5'hc == _T_76[4:0] ? io_in_12_Im : _GEN_716; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_718 = 5'hd == _T_76[4:0] ? io_in_13_Im : _GEN_717; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_719 = 5'he == _T_76[4:0] ? io_in_14_Im : _GEN_718; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_720 = 5'hf == _T_76[4:0] ? io_in_15_Im : _GEN_719; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_721 = 5'h10 == _T_76[4:0] ? io_in_16_Im : _GEN_720; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_722 = 5'h11 == _T_76[4:0] ? io_in_17_Im : _GEN_721; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_723 = 5'h12 == _T_76[4:0] ? io_in_18_Im : _GEN_722; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_724 = 5'h13 == _T_76[4:0] ? io_in_19_Im : _GEN_723; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_725 = 5'h14 == _T_76[4:0] ? io_in_20_Im : _GEN_724; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_726 = 5'h15 == _T_76[4:0] ? io_in_21_Im : _GEN_725; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_727 = 5'h16 == _T_76[4:0] ? io_in_22_Im : _GEN_726; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_728 = 5'h17 == _T_76[4:0] ? io_in_23_Im : _GEN_727; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_729 = 5'h18 == _T_76[4:0] ? io_in_24_Im : _GEN_728; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_730 = 5'h19 == _T_76[4:0] ? io_in_25_Im : _GEN_729; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_733 = 5'h1 == _T_76[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_734 = 5'h2 == _T_76[4:0] ? io_in_2_Re : _GEN_733; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_735 = 5'h3 == _T_76[4:0] ? io_in_3_Re : _GEN_734; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_736 = 5'h4 == _T_76[4:0] ? io_in_4_Re : _GEN_735; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_737 = 5'h5 == _T_76[4:0] ? io_in_5_Re : _GEN_736; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_738 = 5'h6 == _T_76[4:0] ? io_in_6_Re : _GEN_737; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_739 = 5'h7 == _T_76[4:0] ? io_in_7_Re : _GEN_738; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_740 = 5'h8 == _T_76[4:0] ? io_in_8_Re : _GEN_739; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_741 = 5'h9 == _T_76[4:0] ? io_in_9_Re : _GEN_740; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_742 = 5'ha == _T_76[4:0] ? io_in_10_Re : _GEN_741; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_743 = 5'hb == _T_76[4:0] ? io_in_11_Re : _GEN_742; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_744 = 5'hc == _T_76[4:0] ? io_in_12_Re : _GEN_743; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_745 = 5'hd == _T_76[4:0] ? io_in_13_Re : _GEN_744; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_746 = 5'he == _T_76[4:0] ? io_in_14_Re : _GEN_745; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_747 = 5'hf == _T_76[4:0] ? io_in_15_Re : _GEN_746; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_748 = 5'h10 == _T_76[4:0] ? io_in_16_Re : _GEN_747; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_749 = 5'h11 == _T_76[4:0] ? io_in_17_Re : _GEN_748; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_750 = 5'h12 == _T_76[4:0] ? io_in_18_Re : _GEN_749; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_751 = 5'h13 == _T_76[4:0] ? io_in_19_Re : _GEN_750; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_752 = 5'h14 == _T_76[4:0] ? io_in_20_Re : _GEN_751; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_753 = 5'h15 == _T_76[4:0] ? io_in_21_Re : _GEN_752; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_754 = 5'h16 == _T_76[4:0] ? io_in_22_Re : _GEN_753; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_755 = 5'h17 == _T_76[4:0] ? io_in_23_Re : _GEN_754; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_756 = 5'h18 == _T_76[4:0] ? io_in_24_Re : _GEN_755; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_757 = 5'h19 == _T_76[4:0] ? io_in_25_Re : _GEN_756; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_88 = _T_2 + 37'h7; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_769 = 5'ha == _T_88[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_770 = 5'hb == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_769; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_771 = 5'hc == _T_88[4:0] ? 32'h3f800000 : _GEN_770; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_772 = 5'hd == _T_88[4:0] ? 32'h3f441b7c : _GEN_771; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_773 = 5'he == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_772; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_774 = 5'hf == _T_88[4:0] ? 32'h3f800000 : _GEN_773; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_775 = 5'h10 == _T_88[4:0] ? 32'h3f441b7c : _GEN_774; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_776 = 5'h11 == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_775; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_777 = 5'h12 == _T_88[4:0] ? 32'h3f800000 : _GEN_776; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_778 = 5'h13 == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_777; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_779 = 5'h14 == _T_88[4:0] ? 32'hbf708fb2 : _GEN_778; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_780 = 5'h15 == _T_88[4:0] ? 32'h3f800000 : _GEN_779; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_781 = 5'h16 == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_780; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_782 = 5'h17 == _T_88[4:0] ? 32'hbf708fb2 : _GEN_781; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_783 = 5'h18 == _T_88[4:0] ? 32'h3f800000 : _GEN_782; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_784 = 5'h19 == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_783; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_796 = 5'ha == _T_88[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_797 = 5'hb == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_796; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_798 = 5'hc == _T_88[4:0] ? 32'h80800000 : _GEN_797; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_799 = 5'hd == _T_88[4:0] ? 32'hbf248dba : _GEN_798; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_800 = 5'he == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_799; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_801 = 5'hf == _T_88[4:0] ? 32'h80800000 : _GEN_800; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_802 = 5'h10 == _T_88[4:0] ? 32'hbf248dba : _GEN_801; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_803 = 5'h11 == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_802; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_804 = 5'h12 == _T_88[4:0] ? 32'h80800000 : _GEN_803; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_805 = 5'h13 == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_804; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_806 = 5'h14 == _T_88[4:0] ? 32'hbeaf1d40 : _GEN_805; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_807 = 5'h15 == _T_88[4:0] ? 32'h80800000 : _GEN_806; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_808 = 5'h16 == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_807; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_809 = 5'h17 == _T_88[4:0] ? 32'hbeaf1d40 : _GEN_808; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_810 = 5'h18 == _T_88[4:0] ? 32'h80800000 : _GEN_809; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_811 = 5'h19 == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_810; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_814 = 5'h1 == _T_88[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_815 = 5'h2 == _T_88[4:0] ? io_in_2_Im : _GEN_814; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_816 = 5'h3 == _T_88[4:0] ? io_in_3_Im : _GEN_815; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_817 = 5'h4 == _T_88[4:0] ? io_in_4_Im : _GEN_816; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_818 = 5'h5 == _T_88[4:0] ? io_in_5_Im : _GEN_817; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_819 = 5'h6 == _T_88[4:0] ? io_in_6_Im : _GEN_818; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_820 = 5'h7 == _T_88[4:0] ? io_in_7_Im : _GEN_819; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_821 = 5'h8 == _T_88[4:0] ? io_in_8_Im : _GEN_820; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_822 = 5'h9 == _T_88[4:0] ? io_in_9_Im : _GEN_821; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_823 = 5'ha == _T_88[4:0] ? io_in_10_Im : _GEN_822; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_824 = 5'hb == _T_88[4:0] ? io_in_11_Im : _GEN_823; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_825 = 5'hc == _T_88[4:0] ? io_in_12_Im : _GEN_824; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_826 = 5'hd == _T_88[4:0] ? io_in_13_Im : _GEN_825; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_827 = 5'he == _T_88[4:0] ? io_in_14_Im : _GEN_826; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_828 = 5'hf == _T_88[4:0] ? io_in_15_Im : _GEN_827; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_829 = 5'h10 == _T_88[4:0] ? io_in_16_Im : _GEN_828; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_830 = 5'h11 == _T_88[4:0] ? io_in_17_Im : _GEN_829; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_831 = 5'h12 == _T_88[4:0] ? io_in_18_Im : _GEN_830; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_832 = 5'h13 == _T_88[4:0] ? io_in_19_Im : _GEN_831; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_833 = 5'h14 == _T_88[4:0] ? io_in_20_Im : _GEN_832; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_834 = 5'h15 == _T_88[4:0] ? io_in_21_Im : _GEN_833; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_835 = 5'h16 == _T_88[4:0] ? io_in_22_Im : _GEN_834; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_836 = 5'h17 == _T_88[4:0] ? io_in_23_Im : _GEN_835; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_837 = 5'h18 == _T_88[4:0] ? io_in_24_Im : _GEN_836; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_838 = 5'h19 == _T_88[4:0] ? io_in_25_Im : _GEN_837; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_841 = 5'h1 == _T_88[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_842 = 5'h2 == _T_88[4:0] ? io_in_2_Re : _GEN_841; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_843 = 5'h3 == _T_88[4:0] ? io_in_3_Re : _GEN_842; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_844 = 5'h4 == _T_88[4:0] ? io_in_4_Re : _GEN_843; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_845 = 5'h5 == _T_88[4:0] ? io_in_5_Re : _GEN_844; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_846 = 5'h6 == _T_88[4:0] ? io_in_6_Re : _GEN_845; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_847 = 5'h7 == _T_88[4:0] ? io_in_7_Re : _GEN_846; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_848 = 5'h8 == _T_88[4:0] ? io_in_8_Re : _GEN_847; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_849 = 5'h9 == _T_88[4:0] ? io_in_9_Re : _GEN_848; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_850 = 5'ha == _T_88[4:0] ? io_in_10_Re : _GEN_849; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_851 = 5'hb == _T_88[4:0] ? io_in_11_Re : _GEN_850; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_852 = 5'hc == _T_88[4:0] ? io_in_12_Re : _GEN_851; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_853 = 5'hd == _T_88[4:0] ? io_in_13_Re : _GEN_852; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_854 = 5'he == _T_88[4:0] ? io_in_14_Re : _GEN_853; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_855 = 5'hf == _T_88[4:0] ? io_in_15_Re : _GEN_854; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_856 = 5'h10 == _T_88[4:0] ? io_in_16_Re : _GEN_855; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_857 = 5'h11 == _T_88[4:0] ? io_in_17_Re : _GEN_856; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_858 = 5'h12 == _T_88[4:0] ? io_in_18_Re : _GEN_857; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_859 = 5'h13 == _T_88[4:0] ? io_in_19_Re : _GEN_858; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_860 = 5'h14 == _T_88[4:0] ? io_in_20_Re : _GEN_859; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_861 = 5'h15 == _T_88[4:0] ? io_in_21_Re : _GEN_860; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_862 = 5'h16 == _T_88[4:0] ? io_in_22_Re : _GEN_861; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_863 = 5'h17 == _T_88[4:0] ? io_in_23_Re : _GEN_862; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_864 = 5'h18 == _T_88[4:0] ? io_in_24_Re : _GEN_863; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_865 = 5'h19 == _T_88[4:0] ? io_in_25_Re : _GEN_864; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_100 = _T_2 + 37'h8; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_877 = 5'ha == _T_100[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_878 = 5'hb == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_877; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_879 = 5'hc == _T_100[4:0] ? 32'h3f800000 : _GEN_878; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_880 = 5'hd == _T_100[4:0] ? 32'h3f441b7c : _GEN_879; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_881 = 5'he == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_880; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_882 = 5'hf == _T_100[4:0] ? 32'h3f800000 : _GEN_881; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_883 = 5'h10 == _T_100[4:0] ? 32'h3f441b7c : _GEN_882; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_884 = 5'h11 == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_883; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_885 = 5'h12 == _T_100[4:0] ? 32'h3f800000 : _GEN_884; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_886 = 5'h13 == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_885; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_887 = 5'h14 == _T_100[4:0] ? 32'hbf708fb2 : _GEN_886; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_888 = 5'h15 == _T_100[4:0] ? 32'h3f800000 : _GEN_887; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_889 = 5'h16 == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_888; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_890 = 5'h17 == _T_100[4:0] ? 32'hbf708fb2 : _GEN_889; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_891 = 5'h18 == _T_100[4:0] ? 32'h3f800000 : _GEN_890; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_892 = 5'h19 == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_891; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_904 = 5'ha == _T_100[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_905 = 5'hb == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_904; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_906 = 5'hc == _T_100[4:0] ? 32'h80800000 : _GEN_905; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_907 = 5'hd == _T_100[4:0] ? 32'hbf248dba : _GEN_906; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_908 = 5'he == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_907; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_909 = 5'hf == _T_100[4:0] ? 32'h80800000 : _GEN_908; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_910 = 5'h10 == _T_100[4:0] ? 32'hbf248dba : _GEN_909; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_911 = 5'h11 == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_910; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_912 = 5'h12 == _T_100[4:0] ? 32'h80800000 : _GEN_911; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_913 = 5'h13 == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_912; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_914 = 5'h14 == _T_100[4:0] ? 32'hbeaf1d40 : _GEN_913; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_915 = 5'h15 == _T_100[4:0] ? 32'h80800000 : _GEN_914; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_916 = 5'h16 == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_915; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_917 = 5'h17 == _T_100[4:0] ? 32'hbeaf1d40 : _GEN_916; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_918 = 5'h18 == _T_100[4:0] ? 32'h80800000 : _GEN_917; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_919 = 5'h19 == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_918; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_922 = 5'h1 == _T_100[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_923 = 5'h2 == _T_100[4:0] ? io_in_2_Im : _GEN_922; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_924 = 5'h3 == _T_100[4:0] ? io_in_3_Im : _GEN_923; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_925 = 5'h4 == _T_100[4:0] ? io_in_4_Im : _GEN_924; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_926 = 5'h5 == _T_100[4:0] ? io_in_5_Im : _GEN_925; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_927 = 5'h6 == _T_100[4:0] ? io_in_6_Im : _GEN_926; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_928 = 5'h7 == _T_100[4:0] ? io_in_7_Im : _GEN_927; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_929 = 5'h8 == _T_100[4:0] ? io_in_8_Im : _GEN_928; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_930 = 5'h9 == _T_100[4:0] ? io_in_9_Im : _GEN_929; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_931 = 5'ha == _T_100[4:0] ? io_in_10_Im : _GEN_930; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_932 = 5'hb == _T_100[4:0] ? io_in_11_Im : _GEN_931; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_933 = 5'hc == _T_100[4:0] ? io_in_12_Im : _GEN_932; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_934 = 5'hd == _T_100[4:0] ? io_in_13_Im : _GEN_933; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_935 = 5'he == _T_100[4:0] ? io_in_14_Im : _GEN_934; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_936 = 5'hf == _T_100[4:0] ? io_in_15_Im : _GEN_935; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_937 = 5'h10 == _T_100[4:0] ? io_in_16_Im : _GEN_936; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_938 = 5'h11 == _T_100[4:0] ? io_in_17_Im : _GEN_937; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_939 = 5'h12 == _T_100[4:0] ? io_in_18_Im : _GEN_938; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_940 = 5'h13 == _T_100[4:0] ? io_in_19_Im : _GEN_939; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_941 = 5'h14 == _T_100[4:0] ? io_in_20_Im : _GEN_940; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_942 = 5'h15 == _T_100[4:0] ? io_in_21_Im : _GEN_941; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_943 = 5'h16 == _T_100[4:0] ? io_in_22_Im : _GEN_942; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_944 = 5'h17 == _T_100[4:0] ? io_in_23_Im : _GEN_943; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_945 = 5'h18 == _T_100[4:0] ? io_in_24_Im : _GEN_944; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_946 = 5'h19 == _T_100[4:0] ? io_in_25_Im : _GEN_945; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_949 = 5'h1 == _T_100[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_950 = 5'h2 == _T_100[4:0] ? io_in_2_Re : _GEN_949; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_951 = 5'h3 == _T_100[4:0] ? io_in_3_Re : _GEN_950; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_952 = 5'h4 == _T_100[4:0] ? io_in_4_Re : _GEN_951; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_953 = 5'h5 == _T_100[4:0] ? io_in_5_Re : _GEN_952; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_954 = 5'h6 == _T_100[4:0] ? io_in_6_Re : _GEN_953; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_955 = 5'h7 == _T_100[4:0] ? io_in_7_Re : _GEN_954; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_956 = 5'h8 == _T_100[4:0] ? io_in_8_Re : _GEN_955; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_957 = 5'h9 == _T_100[4:0] ? io_in_9_Re : _GEN_956; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_958 = 5'ha == _T_100[4:0] ? io_in_10_Re : _GEN_957; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_959 = 5'hb == _T_100[4:0] ? io_in_11_Re : _GEN_958; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_960 = 5'hc == _T_100[4:0] ? io_in_12_Re : _GEN_959; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_961 = 5'hd == _T_100[4:0] ? io_in_13_Re : _GEN_960; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_962 = 5'he == _T_100[4:0] ? io_in_14_Re : _GEN_961; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_963 = 5'hf == _T_100[4:0] ? io_in_15_Re : _GEN_962; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_964 = 5'h10 == _T_100[4:0] ? io_in_16_Re : _GEN_963; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_965 = 5'h11 == _T_100[4:0] ? io_in_17_Re : _GEN_964; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_966 = 5'h12 == _T_100[4:0] ? io_in_18_Re : _GEN_965; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_967 = 5'h13 == _T_100[4:0] ? io_in_19_Re : _GEN_966; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_968 = 5'h14 == _T_100[4:0] ? io_in_20_Re : _GEN_967; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_969 = 5'h15 == _T_100[4:0] ? io_in_21_Re : _GEN_968; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_970 = 5'h16 == _T_100[4:0] ? io_in_22_Re : _GEN_969; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_971 = 5'h17 == _T_100[4:0] ? io_in_23_Re : _GEN_970; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_972 = 5'h18 == _T_100[4:0] ? io_in_24_Re : _GEN_971; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_973 = 5'h19 == _T_100[4:0] ? io_in_25_Re : _GEN_972; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_112 = _T_2 + 37'h9; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_985 = 5'ha == _T_112[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_986 = 5'hb == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_985; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_987 = 5'hc == _T_112[4:0] ? 32'h3f800000 : _GEN_986; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_988 = 5'hd == _T_112[4:0] ? 32'h3f441b7c : _GEN_987; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_989 = 5'he == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_988; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_990 = 5'hf == _T_112[4:0] ? 32'h3f800000 : _GEN_989; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_991 = 5'h10 == _T_112[4:0] ? 32'h3f441b7c : _GEN_990; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_992 = 5'h11 == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_991; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_993 = 5'h12 == _T_112[4:0] ? 32'h3f800000 : _GEN_992; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_994 = 5'h13 == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_993; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_995 = 5'h14 == _T_112[4:0] ? 32'hbf708fb2 : _GEN_994; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_996 = 5'h15 == _T_112[4:0] ? 32'h3f800000 : _GEN_995; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_997 = 5'h16 == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_996; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_998 = 5'h17 == _T_112[4:0] ? 32'hbf708fb2 : _GEN_997; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_999 = 5'h18 == _T_112[4:0] ? 32'h3f800000 : _GEN_998; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1000 = 5'h19 == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_999; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1012 = 5'ha == _T_112[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1013 = 5'hb == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1012; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1014 = 5'hc == _T_112[4:0] ? 32'h80800000 : _GEN_1013; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1015 = 5'hd == _T_112[4:0] ? 32'hbf248dba : _GEN_1014; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1016 = 5'he == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1015; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1017 = 5'hf == _T_112[4:0] ? 32'h80800000 : _GEN_1016; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1018 = 5'h10 == _T_112[4:0] ? 32'hbf248dba : _GEN_1017; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1019 = 5'h11 == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1018; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1020 = 5'h12 == _T_112[4:0] ? 32'h80800000 : _GEN_1019; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1021 = 5'h13 == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1020; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1022 = 5'h14 == _T_112[4:0] ? 32'hbeaf1d40 : _GEN_1021; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1023 = 5'h15 == _T_112[4:0] ? 32'h80800000 : _GEN_1022; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1024 = 5'h16 == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1023; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1025 = 5'h17 == _T_112[4:0] ? 32'hbeaf1d40 : _GEN_1024; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1026 = 5'h18 == _T_112[4:0] ? 32'h80800000 : _GEN_1025; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1027 = 5'h19 == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1026; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1030 = 5'h1 == _T_112[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1031 = 5'h2 == _T_112[4:0] ? io_in_2_Im : _GEN_1030; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1032 = 5'h3 == _T_112[4:0] ? io_in_3_Im : _GEN_1031; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1033 = 5'h4 == _T_112[4:0] ? io_in_4_Im : _GEN_1032; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1034 = 5'h5 == _T_112[4:0] ? io_in_5_Im : _GEN_1033; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1035 = 5'h6 == _T_112[4:0] ? io_in_6_Im : _GEN_1034; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1036 = 5'h7 == _T_112[4:0] ? io_in_7_Im : _GEN_1035; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1037 = 5'h8 == _T_112[4:0] ? io_in_8_Im : _GEN_1036; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1038 = 5'h9 == _T_112[4:0] ? io_in_9_Im : _GEN_1037; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1039 = 5'ha == _T_112[4:0] ? io_in_10_Im : _GEN_1038; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1040 = 5'hb == _T_112[4:0] ? io_in_11_Im : _GEN_1039; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1041 = 5'hc == _T_112[4:0] ? io_in_12_Im : _GEN_1040; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1042 = 5'hd == _T_112[4:0] ? io_in_13_Im : _GEN_1041; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1043 = 5'he == _T_112[4:0] ? io_in_14_Im : _GEN_1042; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1044 = 5'hf == _T_112[4:0] ? io_in_15_Im : _GEN_1043; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1045 = 5'h10 == _T_112[4:0] ? io_in_16_Im : _GEN_1044; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1046 = 5'h11 == _T_112[4:0] ? io_in_17_Im : _GEN_1045; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1047 = 5'h12 == _T_112[4:0] ? io_in_18_Im : _GEN_1046; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1048 = 5'h13 == _T_112[4:0] ? io_in_19_Im : _GEN_1047; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1049 = 5'h14 == _T_112[4:0] ? io_in_20_Im : _GEN_1048; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1050 = 5'h15 == _T_112[4:0] ? io_in_21_Im : _GEN_1049; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1051 = 5'h16 == _T_112[4:0] ? io_in_22_Im : _GEN_1050; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1052 = 5'h17 == _T_112[4:0] ? io_in_23_Im : _GEN_1051; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1053 = 5'h18 == _T_112[4:0] ? io_in_24_Im : _GEN_1052; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1054 = 5'h19 == _T_112[4:0] ? io_in_25_Im : _GEN_1053; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1057 = 5'h1 == _T_112[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1058 = 5'h2 == _T_112[4:0] ? io_in_2_Re : _GEN_1057; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1059 = 5'h3 == _T_112[4:0] ? io_in_3_Re : _GEN_1058; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1060 = 5'h4 == _T_112[4:0] ? io_in_4_Re : _GEN_1059; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1061 = 5'h5 == _T_112[4:0] ? io_in_5_Re : _GEN_1060; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1062 = 5'h6 == _T_112[4:0] ? io_in_6_Re : _GEN_1061; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1063 = 5'h7 == _T_112[4:0] ? io_in_7_Re : _GEN_1062; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1064 = 5'h8 == _T_112[4:0] ? io_in_8_Re : _GEN_1063; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1065 = 5'h9 == _T_112[4:0] ? io_in_9_Re : _GEN_1064; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1066 = 5'ha == _T_112[4:0] ? io_in_10_Re : _GEN_1065; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1067 = 5'hb == _T_112[4:0] ? io_in_11_Re : _GEN_1066; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1068 = 5'hc == _T_112[4:0] ? io_in_12_Re : _GEN_1067; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1069 = 5'hd == _T_112[4:0] ? io_in_13_Re : _GEN_1068; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1070 = 5'he == _T_112[4:0] ? io_in_14_Re : _GEN_1069; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1071 = 5'hf == _T_112[4:0] ? io_in_15_Re : _GEN_1070; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1072 = 5'h10 == _T_112[4:0] ? io_in_16_Re : _GEN_1071; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1073 = 5'h11 == _T_112[4:0] ? io_in_17_Re : _GEN_1072; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1074 = 5'h12 == _T_112[4:0] ? io_in_18_Re : _GEN_1073; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1075 = 5'h13 == _T_112[4:0] ? io_in_19_Re : _GEN_1074; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1076 = 5'h14 == _T_112[4:0] ? io_in_20_Re : _GEN_1075; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1077 = 5'h15 == _T_112[4:0] ? io_in_21_Re : _GEN_1076; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1078 = 5'h16 == _T_112[4:0] ? io_in_22_Re : _GEN_1077; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1079 = 5'h17 == _T_112[4:0] ? io_in_23_Re : _GEN_1078; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1080 = 5'h18 == _T_112[4:0] ? io_in_24_Re : _GEN_1079; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1081 = 5'h19 == _T_112[4:0] ? io_in_25_Re : _GEN_1080; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_124 = _T_2 + 37'ha; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1093 = 5'ha == _T_124[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1094 = 5'hb == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1093; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1095 = 5'hc == _T_124[4:0] ? 32'h3f800000 : _GEN_1094; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1096 = 5'hd == _T_124[4:0] ? 32'h3f441b7c : _GEN_1095; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1097 = 5'he == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1096; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1098 = 5'hf == _T_124[4:0] ? 32'h3f800000 : _GEN_1097; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1099 = 5'h10 == _T_124[4:0] ? 32'h3f441b7c : _GEN_1098; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1100 = 5'h11 == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1099; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1101 = 5'h12 == _T_124[4:0] ? 32'h3f800000 : _GEN_1100; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1102 = 5'h13 == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1101; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1103 = 5'h14 == _T_124[4:0] ? 32'hbf708fb2 : _GEN_1102; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1104 = 5'h15 == _T_124[4:0] ? 32'h3f800000 : _GEN_1103; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1105 = 5'h16 == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1104; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1106 = 5'h17 == _T_124[4:0] ? 32'hbf708fb2 : _GEN_1105; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1107 = 5'h18 == _T_124[4:0] ? 32'h3f800000 : _GEN_1106; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1108 = 5'h19 == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1107; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1120 = 5'ha == _T_124[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1121 = 5'hb == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1120; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1122 = 5'hc == _T_124[4:0] ? 32'h80800000 : _GEN_1121; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1123 = 5'hd == _T_124[4:0] ? 32'hbf248dba : _GEN_1122; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1124 = 5'he == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1123; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1125 = 5'hf == _T_124[4:0] ? 32'h80800000 : _GEN_1124; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1126 = 5'h10 == _T_124[4:0] ? 32'hbf248dba : _GEN_1125; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1127 = 5'h11 == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1126; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1128 = 5'h12 == _T_124[4:0] ? 32'h80800000 : _GEN_1127; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1129 = 5'h13 == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1128; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1130 = 5'h14 == _T_124[4:0] ? 32'hbeaf1d40 : _GEN_1129; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1131 = 5'h15 == _T_124[4:0] ? 32'h80800000 : _GEN_1130; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1132 = 5'h16 == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1131; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1133 = 5'h17 == _T_124[4:0] ? 32'hbeaf1d40 : _GEN_1132; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1134 = 5'h18 == _T_124[4:0] ? 32'h80800000 : _GEN_1133; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1135 = 5'h19 == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1134; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1138 = 5'h1 == _T_124[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1139 = 5'h2 == _T_124[4:0] ? io_in_2_Im : _GEN_1138; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1140 = 5'h3 == _T_124[4:0] ? io_in_3_Im : _GEN_1139; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1141 = 5'h4 == _T_124[4:0] ? io_in_4_Im : _GEN_1140; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1142 = 5'h5 == _T_124[4:0] ? io_in_5_Im : _GEN_1141; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1143 = 5'h6 == _T_124[4:0] ? io_in_6_Im : _GEN_1142; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1144 = 5'h7 == _T_124[4:0] ? io_in_7_Im : _GEN_1143; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1145 = 5'h8 == _T_124[4:0] ? io_in_8_Im : _GEN_1144; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1146 = 5'h9 == _T_124[4:0] ? io_in_9_Im : _GEN_1145; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1147 = 5'ha == _T_124[4:0] ? io_in_10_Im : _GEN_1146; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1148 = 5'hb == _T_124[4:0] ? io_in_11_Im : _GEN_1147; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1149 = 5'hc == _T_124[4:0] ? io_in_12_Im : _GEN_1148; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1150 = 5'hd == _T_124[4:0] ? io_in_13_Im : _GEN_1149; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1151 = 5'he == _T_124[4:0] ? io_in_14_Im : _GEN_1150; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1152 = 5'hf == _T_124[4:0] ? io_in_15_Im : _GEN_1151; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1153 = 5'h10 == _T_124[4:0] ? io_in_16_Im : _GEN_1152; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1154 = 5'h11 == _T_124[4:0] ? io_in_17_Im : _GEN_1153; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1155 = 5'h12 == _T_124[4:0] ? io_in_18_Im : _GEN_1154; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1156 = 5'h13 == _T_124[4:0] ? io_in_19_Im : _GEN_1155; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1157 = 5'h14 == _T_124[4:0] ? io_in_20_Im : _GEN_1156; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1158 = 5'h15 == _T_124[4:0] ? io_in_21_Im : _GEN_1157; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1159 = 5'h16 == _T_124[4:0] ? io_in_22_Im : _GEN_1158; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1160 = 5'h17 == _T_124[4:0] ? io_in_23_Im : _GEN_1159; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1161 = 5'h18 == _T_124[4:0] ? io_in_24_Im : _GEN_1160; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1162 = 5'h19 == _T_124[4:0] ? io_in_25_Im : _GEN_1161; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1165 = 5'h1 == _T_124[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1166 = 5'h2 == _T_124[4:0] ? io_in_2_Re : _GEN_1165; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1167 = 5'h3 == _T_124[4:0] ? io_in_3_Re : _GEN_1166; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1168 = 5'h4 == _T_124[4:0] ? io_in_4_Re : _GEN_1167; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1169 = 5'h5 == _T_124[4:0] ? io_in_5_Re : _GEN_1168; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1170 = 5'h6 == _T_124[4:0] ? io_in_6_Re : _GEN_1169; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1171 = 5'h7 == _T_124[4:0] ? io_in_7_Re : _GEN_1170; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1172 = 5'h8 == _T_124[4:0] ? io_in_8_Re : _GEN_1171; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1173 = 5'h9 == _T_124[4:0] ? io_in_9_Re : _GEN_1172; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1174 = 5'ha == _T_124[4:0] ? io_in_10_Re : _GEN_1173; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1175 = 5'hb == _T_124[4:0] ? io_in_11_Re : _GEN_1174; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1176 = 5'hc == _T_124[4:0] ? io_in_12_Re : _GEN_1175; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1177 = 5'hd == _T_124[4:0] ? io_in_13_Re : _GEN_1176; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1178 = 5'he == _T_124[4:0] ? io_in_14_Re : _GEN_1177; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1179 = 5'hf == _T_124[4:0] ? io_in_15_Re : _GEN_1178; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1180 = 5'h10 == _T_124[4:0] ? io_in_16_Re : _GEN_1179; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1181 = 5'h11 == _T_124[4:0] ? io_in_17_Re : _GEN_1180; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1182 = 5'h12 == _T_124[4:0] ? io_in_18_Re : _GEN_1181; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1183 = 5'h13 == _T_124[4:0] ? io_in_19_Re : _GEN_1182; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1184 = 5'h14 == _T_124[4:0] ? io_in_20_Re : _GEN_1183; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1185 = 5'h15 == _T_124[4:0] ? io_in_21_Re : _GEN_1184; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1186 = 5'h16 == _T_124[4:0] ? io_in_22_Re : _GEN_1185; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1187 = 5'h17 == _T_124[4:0] ? io_in_23_Re : _GEN_1186; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1188 = 5'h18 == _T_124[4:0] ? io_in_24_Re : _GEN_1187; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1189 = 5'h19 == _T_124[4:0] ? io_in_25_Re : _GEN_1188; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_136 = _T_2 + 37'hb; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1201 = 5'ha == _T_136[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1202 = 5'hb == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1201; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1203 = 5'hc == _T_136[4:0] ? 32'h3f800000 : _GEN_1202; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1204 = 5'hd == _T_136[4:0] ? 32'h3f441b7c : _GEN_1203; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1205 = 5'he == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1204; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1206 = 5'hf == _T_136[4:0] ? 32'h3f800000 : _GEN_1205; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1207 = 5'h10 == _T_136[4:0] ? 32'h3f441b7c : _GEN_1206; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1208 = 5'h11 == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1207; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1209 = 5'h12 == _T_136[4:0] ? 32'h3f800000 : _GEN_1208; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1210 = 5'h13 == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1209; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1211 = 5'h14 == _T_136[4:0] ? 32'hbf708fb2 : _GEN_1210; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1212 = 5'h15 == _T_136[4:0] ? 32'h3f800000 : _GEN_1211; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1213 = 5'h16 == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1212; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1214 = 5'h17 == _T_136[4:0] ? 32'hbf708fb2 : _GEN_1213; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1215 = 5'h18 == _T_136[4:0] ? 32'h3f800000 : _GEN_1214; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1216 = 5'h19 == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1215; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1228 = 5'ha == _T_136[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1229 = 5'hb == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1228; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1230 = 5'hc == _T_136[4:0] ? 32'h80800000 : _GEN_1229; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1231 = 5'hd == _T_136[4:0] ? 32'hbf248dba : _GEN_1230; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1232 = 5'he == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1231; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1233 = 5'hf == _T_136[4:0] ? 32'h80800000 : _GEN_1232; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1234 = 5'h10 == _T_136[4:0] ? 32'hbf248dba : _GEN_1233; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1235 = 5'h11 == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1234; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1236 = 5'h12 == _T_136[4:0] ? 32'h80800000 : _GEN_1235; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1237 = 5'h13 == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1236; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1238 = 5'h14 == _T_136[4:0] ? 32'hbeaf1d40 : _GEN_1237; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1239 = 5'h15 == _T_136[4:0] ? 32'h80800000 : _GEN_1238; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1240 = 5'h16 == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1239; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1241 = 5'h17 == _T_136[4:0] ? 32'hbeaf1d40 : _GEN_1240; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1242 = 5'h18 == _T_136[4:0] ? 32'h80800000 : _GEN_1241; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1243 = 5'h19 == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1242; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1246 = 5'h1 == _T_136[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1247 = 5'h2 == _T_136[4:0] ? io_in_2_Im : _GEN_1246; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1248 = 5'h3 == _T_136[4:0] ? io_in_3_Im : _GEN_1247; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1249 = 5'h4 == _T_136[4:0] ? io_in_4_Im : _GEN_1248; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1250 = 5'h5 == _T_136[4:0] ? io_in_5_Im : _GEN_1249; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1251 = 5'h6 == _T_136[4:0] ? io_in_6_Im : _GEN_1250; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1252 = 5'h7 == _T_136[4:0] ? io_in_7_Im : _GEN_1251; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1253 = 5'h8 == _T_136[4:0] ? io_in_8_Im : _GEN_1252; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1254 = 5'h9 == _T_136[4:0] ? io_in_9_Im : _GEN_1253; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1255 = 5'ha == _T_136[4:0] ? io_in_10_Im : _GEN_1254; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1256 = 5'hb == _T_136[4:0] ? io_in_11_Im : _GEN_1255; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1257 = 5'hc == _T_136[4:0] ? io_in_12_Im : _GEN_1256; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1258 = 5'hd == _T_136[4:0] ? io_in_13_Im : _GEN_1257; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1259 = 5'he == _T_136[4:0] ? io_in_14_Im : _GEN_1258; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1260 = 5'hf == _T_136[4:0] ? io_in_15_Im : _GEN_1259; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1261 = 5'h10 == _T_136[4:0] ? io_in_16_Im : _GEN_1260; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1262 = 5'h11 == _T_136[4:0] ? io_in_17_Im : _GEN_1261; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1263 = 5'h12 == _T_136[4:0] ? io_in_18_Im : _GEN_1262; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1264 = 5'h13 == _T_136[4:0] ? io_in_19_Im : _GEN_1263; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1265 = 5'h14 == _T_136[4:0] ? io_in_20_Im : _GEN_1264; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1266 = 5'h15 == _T_136[4:0] ? io_in_21_Im : _GEN_1265; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1267 = 5'h16 == _T_136[4:0] ? io_in_22_Im : _GEN_1266; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1268 = 5'h17 == _T_136[4:0] ? io_in_23_Im : _GEN_1267; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1269 = 5'h18 == _T_136[4:0] ? io_in_24_Im : _GEN_1268; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1270 = 5'h19 == _T_136[4:0] ? io_in_25_Im : _GEN_1269; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1273 = 5'h1 == _T_136[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1274 = 5'h2 == _T_136[4:0] ? io_in_2_Re : _GEN_1273; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1275 = 5'h3 == _T_136[4:0] ? io_in_3_Re : _GEN_1274; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1276 = 5'h4 == _T_136[4:0] ? io_in_4_Re : _GEN_1275; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1277 = 5'h5 == _T_136[4:0] ? io_in_5_Re : _GEN_1276; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1278 = 5'h6 == _T_136[4:0] ? io_in_6_Re : _GEN_1277; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1279 = 5'h7 == _T_136[4:0] ? io_in_7_Re : _GEN_1278; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1280 = 5'h8 == _T_136[4:0] ? io_in_8_Re : _GEN_1279; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1281 = 5'h9 == _T_136[4:0] ? io_in_9_Re : _GEN_1280; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1282 = 5'ha == _T_136[4:0] ? io_in_10_Re : _GEN_1281; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1283 = 5'hb == _T_136[4:0] ? io_in_11_Re : _GEN_1282; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1284 = 5'hc == _T_136[4:0] ? io_in_12_Re : _GEN_1283; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1285 = 5'hd == _T_136[4:0] ? io_in_13_Re : _GEN_1284; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1286 = 5'he == _T_136[4:0] ? io_in_14_Re : _GEN_1285; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1287 = 5'hf == _T_136[4:0] ? io_in_15_Re : _GEN_1286; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1288 = 5'h10 == _T_136[4:0] ? io_in_16_Re : _GEN_1287; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1289 = 5'h11 == _T_136[4:0] ? io_in_17_Re : _GEN_1288; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1290 = 5'h12 == _T_136[4:0] ? io_in_18_Re : _GEN_1289; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1291 = 5'h13 == _T_136[4:0] ? io_in_19_Re : _GEN_1290; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1292 = 5'h14 == _T_136[4:0] ? io_in_20_Re : _GEN_1291; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1293 = 5'h15 == _T_136[4:0] ? io_in_21_Re : _GEN_1292; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1294 = 5'h16 == _T_136[4:0] ? io_in_22_Re : _GEN_1293; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1295 = 5'h17 == _T_136[4:0] ? io_in_23_Re : _GEN_1294; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1296 = 5'h18 == _T_136[4:0] ? io_in_24_Re : _GEN_1295; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1297 = 5'h19 == _T_136[4:0] ? io_in_25_Re : _GEN_1296; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_148 = _T_2 + 37'hc; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1309 = 5'ha == _T_148[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1310 = 5'hb == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1309; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1311 = 5'hc == _T_148[4:0] ? 32'h3f800000 : _GEN_1310; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1312 = 5'hd == _T_148[4:0] ? 32'h3f441b7c : _GEN_1311; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1313 = 5'he == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1312; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1314 = 5'hf == _T_148[4:0] ? 32'h3f800000 : _GEN_1313; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1315 = 5'h10 == _T_148[4:0] ? 32'h3f441b7c : _GEN_1314; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1316 = 5'h11 == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1315; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1317 = 5'h12 == _T_148[4:0] ? 32'h3f800000 : _GEN_1316; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1318 = 5'h13 == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1317; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1319 = 5'h14 == _T_148[4:0] ? 32'hbf708fb2 : _GEN_1318; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1320 = 5'h15 == _T_148[4:0] ? 32'h3f800000 : _GEN_1319; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1321 = 5'h16 == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1320; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1322 = 5'h17 == _T_148[4:0] ? 32'hbf708fb2 : _GEN_1321; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1323 = 5'h18 == _T_148[4:0] ? 32'h3f800000 : _GEN_1322; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1324 = 5'h19 == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1323; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1336 = 5'ha == _T_148[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1337 = 5'hb == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1336; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1338 = 5'hc == _T_148[4:0] ? 32'h80800000 : _GEN_1337; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1339 = 5'hd == _T_148[4:0] ? 32'hbf248dba : _GEN_1338; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1340 = 5'he == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1339; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1341 = 5'hf == _T_148[4:0] ? 32'h80800000 : _GEN_1340; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1342 = 5'h10 == _T_148[4:0] ? 32'hbf248dba : _GEN_1341; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1343 = 5'h11 == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1342; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1344 = 5'h12 == _T_148[4:0] ? 32'h80800000 : _GEN_1343; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1345 = 5'h13 == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1344; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1346 = 5'h14 == _T_148[4:0] ? 32'hbeaf1d40 : _GEN_1345; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1347 = 5'h15 == _T_148[4:0] ? 32'h80800000 : _GEN_1346; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1348 = 5'h16 == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1347; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1349 = 5'h17 == _T_148[4:0] ? 32'hbeaf1d40 : _GEN_1348; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1350 = 5'h18 == _T_148[4:0] ? 32'h80800000 : _GEN_1349; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1351 = 5'h19 == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1350; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1354 = 5'h1 == _T_148[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1355 = 5'h2 == _T_148[4:0] ? io_in_2_Im : _GEN_1354; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1356 = 5'h3 == _T_148[4:0] ? io_in_3_Im : _GEN_1355; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1357 = 5'h4 == _T_148[4:0] ? io_in_4_Im : _GEN_1356; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1358 = 5'h5 == _T_148[4:0] ? io_in_5_Im : _GEN_1357; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1359 = 5'h6 == _T_148[4:0] ? io_in_6_Im : _GEN_1358; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1360 = 5'h7 == _T_148[4:0] ? io_in_7_Im : _GEN_1359; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1361 = 5'h8 == _T_148[4:0] ? io_in_8_Im : _GEN_1360; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1362 = 5'h9 == _T_148[4:0] ? io_in_9_Im : _GEN_1361; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1363 = 5'ha == _T_148[4:0] ? io_in_10_Im : _GEN_1362; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1364 = 5'hb == _T_148[4:0] ? io_in_11_Im : _GEN_1363; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1365 = 5'hc == _T_148[4:0] ? io_in_12_Im : _GEN_1364; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1366 = 5'hd == _T_148[4:0] ? io_in_13_Im : _GEN_1365; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1367 = 5'he == _T_148[4:0] ? io_in_14_Im : _GEN_1366; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1368 = 5'hf == _T_148[4:0] ? io_in_15_Im : _GEN_1367; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1369 = 5'h10 == _T_148[4:0] ? io_in_16_Im : _GEN_1368; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1370 = 5'h11 == _T_148[4:0] ? io_in_17_Im : _GEN_1369; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1371 = 5'h12 == _T_148[4:0] ? io_in_18_Im : _GEN_1370; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1372 = 5'h13 == _T_148[4:0] ? io_in_19_Im : _GEN_1371; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1373 = 5'h14 == _T_148[4:0] ? io_in_20_Im : _GEN_1372; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1374 = 5'h15 == _T_148[4:0] ? io_in_21_Im : _GEN_1373; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1375 = 5'h16 == _T_148[4:0] ? io_in_22_Im : _GEN_1374; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1376 = 5'h17 == _T_148[4:0] ? io_in_23_Im : _GEN_1375; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1377 = 5'h18 == _T_148[4:0] ? io_in_24_Im : _GEN_1376; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1378 = 5'h19 == _T_148[4:0] ? io_in_25_Im : _GEN_1377; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1381 = 5'h1 == _T_148[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1382 = 5'h2 == _T_148[4:0] ? io_in_2_Re : _GEN_1381; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1383 = 5'h3 == _T_148[4:0] ? io_in_3_Re : _GEN_1382; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1384 = 5'h4 == _T_148[4:0] ? io_in_4_Re : _GEN_1383; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1385 = 5'h5 == _T_148[4:0] ? io_in_5_Re : _GEN_1384; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1386 = 5'h6 == _T_148[4:0] ? io_in_6_Re : _GEN_1385; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1387 = 5'h7 == _T_148[4:0] ? io_in_7_Re : _GEN_1386; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1388 = 5'h8 == _T_148[4:0] ? io_in_8_Re : _GEN_1387; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1389 = 5'h9 == _T_148[4:0] ? io_in_9_Re : _GEN_1388; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1390 = 5'ha == _T_148[4:0] ? io_in_10_Re : _GEN_1389; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1391 = 5'hb == _T_148[4:0] ? io_in_11_Re : _GEN_1390; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1392 = 5'hc == _T_148[4:0] ? io_in_12_Re : _GEN_1391; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1393 = 5'hd == _T_148[4:0] ? io_in_13_Re : _GEN_1392; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1394 = 5'he == _T_148[4:0] ? io_in_14_Re : _GEN_1393; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1395 = 5'hf == _T_148[4:0] ? io_in_15_Re : _GEN_1394; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1396 = 5'h10 == _T_148[4:0] ? io_in_16_Re : _GEN_1395; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1397 = 5'h11 == _T_148[4:0] ? io_in_17_Re : _GEN_1396; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1398 = 5'h12 == _T_148[4:0] ? io_in_18_Re : _GEN_1397; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1399 = 5'h13 == _T_148[4:0] ? io_in_19_Re : _GEN_1398; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1400 = 5'h14 == _T_148[4:0] ? io_in_20_Re : _GEN_1399; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1401 = 5'h15 == _T_148[4:0] ? io_in_21_Re : _GEN_1400; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1402 = 5'h16 == _T_148[4:0] ? io_in_22_Re : _GEN_1401; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1403 = 5'h17 == _T_148[4:0] ? io_in_23_Re : _GEN_1402; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1404 = 5'h18 == _T_148[4:0] ? io_in_24_Re : _GEN_1403; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1405 = 5'h19 == _T_148[4:0] ? io_in_25_Re : _GEN_1404; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_160 = _T_2 + 37'hd; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1417 = 5'ha == _T_160[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1418 = 5'hb == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1417; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1419 = 5'hc == _T_160[4:0] ? 32'h3f800000 : _GEN_1418; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1420 = 5'hd == _T_160[4:0] ? 32'h3f441b7c : _GEN_1419; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1421 = 5'he == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1420; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1422 = 5'hf == _T_160[4:0] ? 32'h3f800000 : _GEN_1421; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1423 = 5'h10 == _T_160[4:0] ? 32'h3f441b7c : _GEN_1422; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1424 = 5'h11 == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1423; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1425 = 5'h12 == _T_160[4:0] ? 32'h3f800000 : _GEN_1424; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1426 = 5'h13 == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1425; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1427 = 5'h14 == _T_160[4:0] ? 32'hbf708fb2 : _GEN_1426; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1428 = 5'h15 == _T_160[4:0] ? 32'h3f800000 : _GEN_1427; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1429 = 5'h16 == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1428; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1430 = 5'h17 == _T_160[4:0] ? 32'hbf708fb2 : _GEN_1429; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1431 = 5'h18 == _T_160[4:0] ? 32'h3f800000 : _GEN_1430; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1432 = 5'h19 == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1431; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1444 = 5'ha == _T_160[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1445 = 5'hb == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1444; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1446 = 5'hc == _T_160[4:0] ? 32'h80800000 : _GEN_1445; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1447 = 5'hd == _T_160[4:0] ? 32'hbf248dba : _GEN_1446; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1448 = 5'he == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1447; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1449 = 5'hf == _T_160[4:0] ? 32'h80800000 : _GEN_1448; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1450 = 5'h10 == _T_160[4:0] ? 32'hbf248dba : _GEN_1449; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1451 = 5'h11 == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1450; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1452 = 5'h12 == _T_160[4:0] ? 32'h80800000 : _GEN_1451; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1453 = 5'h13 == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1452; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1454 = 5'h14 == _T_160[4:0] ? 32'hbeaf1d40 : _GEN_1453; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1455 = 5'h15 == _T_160[4:0] ? 32'h80800000 : _GEN_1454; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1456 = 5'h16 == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1455; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1457 = 5'h17 == _T_160[4:0] ? 32'hbeaf1d40 : _GEN_1456; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1458 = 5'h18 == _T_160[4:0] ? 32'h80800000 : _GEN_1457; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1459 = 5'h19 == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1458; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1462 = 5'h1 == _T_160[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1463 = 5'h2 == _T_160[4:0] ? io_in_2_Im : _GEN_1462; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1464 = 5'h3 == _T_160[4:0] ? io_in_3_Im : _GEN_1463; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1465 = 5'h4 == _T_160[4:0] ? io_in_4_Im : _GEN_1464; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1466 = 5'h5 == _T_160[4:0] ? io_in_5_Im : _GEN_1465; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1467 = 5'h6 == _T_160[4:0] ? io_in_6_Im : _GEN_1466; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1468 = 5'h7 == _T_160[4:0] ? io_in_7_Im : _GEN_1467; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1469 = 5'h8 == _T_160[4:0] ? io_in_8_Im : _GEN_1468; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1470 = 5'h9 == _T_160[4:0] ? io_in_9_Im : _GEN_1469; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1471 = 5'ha == _T_160[4:0] ? io_in_10_Im : _GEN_1470; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1472 = 5'hb == _T_160[4:0] ? io_in_11_Im : _GEN_1471; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1473 = 5'hc == _T_160[4:0] ? io_in_12_Im : _GEN_1472; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1474 = 5'hd == _T_160[4:0] ? io_in_13_Im : _GEN_1473; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1475 = 5'he == _T_160[4:0] ? io_in_14_Im : _GEN_1474; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1476 = 5'hf == _T_160[4:0] ? io_in_15_Im : _GEN_1475; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1477 = 5'h10 == _T_160[4:0] ? io_in_16_Im : _GEN_1476; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1478 = 5'h11 == _T_160[4:0] ? io_in_17_Im : _GEN_1477; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1479 = 5'h12 == _T_160[4:0] ? io_in_18_Im : _GEN_1478; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1480 = 5'h13 == _T_160[4:0] ? io_in_19_Im : _GEN_1479; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1481 = 5'h14 == _T_160[4:0] ? io_in_20_Im : _GEN_1480; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1482 = 5'h15 == _T_160[4:0] ? io_in_21_Im : _GEN_1481; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1483 = 5'h16 == _T_160[4:0] ? io_in_22_Im : _GEN_1482; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1484 = 5'h17 == _T_160[4:0] ? io_in_23_Im : _GEN_1483; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1485 = 5'h18 == _T_160[4:0] ? io_in_24_Im : _GEN_1484; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1486 = 5'h19 == _T_160[4:0] ? io_in_25_Im : _GEN_1485; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1489 = 5'h1 == _T_160[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1490 = 5'h2 == _T_160[4:0] ? io_in_2_Re : _GEN_1489; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1491 = 5'h3 == _T_160[4:0] ? io_in_3_Re : _GEN_1490; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1492 = 5'h4 == _T_160[4:0] ? io_in_4_Re : _GEN_1491; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1493 = 5'h5 == _T_160[4:0] ? io_in_5_Re : _GEN_1492; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1494 = 5'h6 == _T_160[4:0] ? io_in_6_Re : _GEN_1493; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1495 = 5'h7 == _T_160[4:0] ? io_in_7_Re : _GEN_1494; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1496 = 5'h8 == _T_160[4:0] ? io_in_8_Re : _GEN_1495; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1497 = 5'h9 == _T_160[4:0] ? io_in_9_Re : _GEN_1496; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1498 = 5'ha == _T_160[4:0] ? io_in_10_Re : _GEN_1497; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1499 = 5'hb == _T_160[4:0] ? io_in_11_Re : _GEN_1498; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1500 = 5'hc == _T_160[4:0] ? io_in_12_Re : _GEN_1499; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1501 = 5'hd == _T_160[4:0] ? io_in_13_Re : _GEN_1500; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1502 = 5'he == _T_160[4:0] ? io_in_14_Re : _GEN_1501; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1503 = 5'hf == _T_160[4:0] ? io_in_15_Re : _GEN_1502; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1504 = 5'h10 == _T_160[4:0] ? io_in_16_Re : _GEN_1503; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1505 = 5'h11 == _T_160[4:0] ? io_in_17_Re : _GEN_1504; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1506 = 5'h12 == _T_160[4:0] ? io_in_18_Re : _GEN_1505; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1507 = 5'h13 == _T_160[4:0] ? io_in_19_Re : _GEN_1506; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1508 = 5'h14 == _T_160[4:0] ? io_in_20_Re : _GEN_1507; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1509 = 5'h15 == _T_160[4:0] ? io_in_21_Re : _GEN_1508; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1510 = 5'h16 == _T_160[4:0] ? io_in_22_Re : _GEN_1509; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1511 = 5'h17 == _T_160[4:0] ? io_in_23_Re : _GEN_1510; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1512 = 5'h18 == _T_160[4:0] ? io_in_24_Re : _GEN_1511; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1513 = 5'h19 == _T_160[4:0] ? io_in_25_Re : _GEN_1512; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_172 = _T_2 + 37'he; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1525 = 5'ha == _T_172[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1526 = 5'hb == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1525; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1527 = 5'hc == _T_172[4:0] ? 32'h3f800000 : _GEN_1526; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1528 = 5'hd == _T_172[4:0] ? 32'h3f441b7c : _GEN_1527; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1529 = 5'he == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1528; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1530 = 5'hf == _T_172[4:0] ? 32'h3f800000 : _GEN_1529; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1531 = 5'h10 == _T_172[4:0] ? 32'h3f441b7c : _GEN_1530; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1532 = 5'h11 == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1531; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1533 = 5'h12 == _T_172[4:0] ? 32'h3f800000 : _GEN_1532; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1534 = 5'h13 == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1533; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1535 = 5'h14 == _T_172[4:0] ? 32'hbf708fb2 : _GEN_1534; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1536 = 5'h15 == _T_172[4:0] ? 32'h3f800000 : _GEN_1535; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1537 = 5'h16 == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1536; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1538 = 5'h17 == _T_172[4:0] ? 32'hbf708fb2 : _GEN_1537; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1539 = 5'h18 == _T_172[4:0] ? 32'h3f800000 : _GEN_1538; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1540 = 5'h19 == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1539; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1552 = 5'ha == _T_172[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1553 = 5'hb == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1552; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1554 = 5'hc == _T_172[4:0] ? 32'h80800000 : _GEN_1553; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1555 = 5'hd == _T_172[4:0] ? 32'hbf248dba : _GEN_1554; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1556 = 5'he == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1555; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1557 = 5'hf == _T_172[4:0] ? 32'h80800000 : _GEN_1556; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1558 = 5'h10 == _T_172[4:0] ? 32'hbf248dba : _GEN_1557; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1559 = 5'h11 == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1558; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1560 = 5'h12 == _T_172[4:0] ? 32'h80800000 : _GEN_1559; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1561 = 5'h13 == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1560; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1562 = 5'h14 == _T_172[4:0] ? 32'hbeaf1d40 : _GEN_1561; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1563 = 5'h15 == _T_172[4:0] ? 32'h80800000 : _GEN_1562; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1564 = 5'h16 == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1563; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1565 = 5'h17 == _T_172[4:0] ? 32'hbeaf1d40 : _GEN_1564; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1566 = 5'h18 == _T_172[4:0] ? 32'h80800000 : _GEN_1565; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1567 = 5'h19 == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1566; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1570 = 5'h1 == _T_172[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1571 = 5'h2 == _T_172[4:0] ? io_in_2_Im : _GEN_1570; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1572 = 5'h3 == _T_172[4:0] ? io_in_3_Im : _GEN_1571; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1573 = 5'h4 == _T_172[4:0] ? io_in_4_Im : _GEN_1572; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1574 = 5'h5 == _T_172[4:0] ? io_in_5_Im : _GEN_1573; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1575 = 5'h6 == _T_172[4:0] ? io_in_6_Im : _GEN_1574; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1576 = 5'h7 == _T_172[4:0] ? io_in_7_Im : _GEN_1575; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1577 = 5'h8 == _T_172[4:0] ? io_in_8_Im : _GEN_1576; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1578 = 5'h9 == _T_172[4:0] ? io_in_9_Im : _GEN_1577; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1579 = 5'ha == _T_172[4:0] ? io_in_10_Im : _GEN_1578; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1580 = 5'hb == _T_172[4:0] ? io_in_11_Im : _GEN_1579; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1581 = 5'hc == _T_172[4:0] ? io_in_12_Im : _GEN_1580; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1582 = 5'hd == _T_172[4:0] ? io_in_13_Im : _GEN_1581; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1583 = 5'he == _T_172[4:0] ? io_in_14_Im : _GEN_1582; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1584 = 5'hf == _T_172[4:0] ? io_in_15_Im : _GEN_1583; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1585 = 5'h10 == _T_172[4:0] ? io_in_16_Im : _GEN_1584; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1586 = 5'h11 == _T_172[4:0] ? io_in_17_Im : _GEN_1585; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1587 = 5'h12 == _T_172[4:0] ? io_in_18_Im : _GEN_1586; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1588 = 5'h13 == _T_172[4:0] ? io_in_19_Im : _GEN_1587; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1589 = 5'h14 == _T_172[4:0] ? io_in_20_Im : _GEN_1588; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1590 = 5'h15 == _T_172[4:0] ? io_in_21_Im : _GEN_1589; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1591 = 5'h16 == _T_172[4:0] ? io_in_22_Im : _GEN_1590; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1592 = 5'h17 == _T_172[4:0] ? io_in_23_Im : _GEN_1591; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1593 = 5'h18 == _T_172[4:0] ? io_in_24_Im : _GEN_1592; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1594 = 5'h19 == _T_172[4:0] ? io_in_25_Im : _GEN_1593; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1597 = 5'h1 == _T_172[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1598 = 5'h2 == _T_172[4:0] ? io_in_2_Re : _GEN_1597; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1599 = 5'h3 == _T_172[4:0] ? io_in_3_Re : _GEN_1598; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1600 = 5'h4 == _T_172[4:0] ? io_in_4_Re : _GEN_1599; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1601 = 5'h5 == _T_172[4:0] ? io_in_5_Re : _GEN_1600; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1602 = 5'h6 == _T_172[4:0] ? io_in_6_Re : _GEN_1601; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1603 = 5'h7 == _T_172[4:0] ? io_in_7_Re : _GEN_1602; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1604 = 5'h8 == _T_172[4:0] ? io_in_8_Re : _GEN_1603; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1605 = 5'h9 == _T_172[4:0] ? io_in_9_Re : _GEN_1604; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1606 = 5'ha == _T_172[4:0] ? io_in_10_Re : _GEN_1605; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1607 = 5'hb == _T_172[4:0] ? io_in_11_Re : _GEN_1606; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1608 = 5'hc == _T_172[4:0] ? io_in_12_Re : _GEN_1607; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1609 = 5'hd == _T_172[4:0] ? io_in_13_Re : _GEN_1608; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1610 = 5'he == _T_172[4:0] ? io_in_14_Re : _GEN_1609; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1611 = 5'hf == _T_172[4:0] ? io_in_15_Re : _GEN_1610; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1612 = 5'h10 == _T_172[4:0] ? io_in_16_Re : _GEN_1611; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1613 = 5'h11 == _T_172[4:0] ? io_in_17_Re : _GEN_1612; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1614 = 5'h12 == _T_172[4:0] ? io_in_18_Re : _GEN_1613; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1615 = 5'h13 == _T_172[4:0] ? io_in_19_Re : _GEN_1614; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1616 = 5'h14 == _T_172[4:0] ? io_in_20_Re : _GEN_1615; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1617 = 5'h15 == _T_172[4:0] ? io_in_21_Re : _GEN_1616; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1618 = 5'h16 == _T_172[4:0] ? io_in_22_Re : _GEN_1617; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1619 = 5'h17 == _T_172[4:0] ? io_in_23_Re : _GEN_1618; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1620 = 5'h18 == _T_172[4:0] ? io_in_24_Re : _GEN_1619; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1621 = 5'h19 == _T_172[4:0] ? io_in_25_Re : _GEN_1620; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_184 = _T_2 + 37'hf; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1633 = 5'ha == _T_184[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1634 = 5'hb == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1633; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1635 = 5'hc == _T_184[4:0] ? 32'h3f800000 : _GEN_1634; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1636 = 5'hd == _T_184[4:0] ? 32'h3f441b7c : _GEN_1635; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1637 = 5'he == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1636; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1638 = 5'hf == _T_184[4:0] ? 32'h3f800000 : _GEN_1637; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1639 = 5'h10 == _T_184[4:0] ? 32'h3f441b7c : _GEN_1638; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1640 = 5'h11 == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1639; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1641 = 5'h12 == _T_184[4:0] ? 32'h3f800000 : _GEN_1640; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1642 = 5'h13 == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1641; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1643 = 5'h14 == _T_184[4:0] ? 32'hbf708fb2 : _GEN_1642; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1644 = 5'h15 == _T_184[4:0] ? 32'h3f800000 : _GEN_1643; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1645 = 5'h16 == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1644; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1646 = 5'h17 == _T_184[4:0] ? 32'hbf708fb2 : _GEN_1645; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1647 = 5'h18 == _T_184[4:0] ? 32'h3f800000 : _GEN_1646; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1648 = 5'h19 == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1647; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1660 = 5'ha == _T_184[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1661 = 5'hb == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1660; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1662 = 5'hc == _T_184[4:0] ? 32'h80800000 : _GEN_1661; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1663 = 5'hd == _T_184[4:0] ? 32'hbf248dba : _GEN_1662; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1664 = 5'he == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1663; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1665 = 5'hf == _T_184[4:0] ? 32'h80800000 : _GEN_1664; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1666 = 5'h10 == _T_184[4:0] ? 32'hbf248dba : _GEN_1665; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1667 = 5'h11 == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1666; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1668 = 5'h12 == _T_184[4:0] ? 32'h80800000 : _GEN_1667; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1669 = 5'h13 == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1668; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1670 = 5'h14 == _T_184[4:0] ? 32'hbeaf1d40 : _GEN_1669; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1671 = 5'h15 == _T_184[4:0] ? 32'h80800000 : _GEN_1670; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1672 = 5'h16 == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1671; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1673 = 5'h17 == _T_184[4:0] ? 32'hbeaf1d40 : _GEN_1672; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1674 = 5'h18 == _T_184[4:0] ? 32'h80800000 : _GEN_1673; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1675 = 5'h19 == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1674; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1678 = 5'h1 == _T_184[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1679 = 5'h2 == _T_184[4:0] ? io_in_2_Im : _GEN_1678; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1680 = 5'h3 == _T_184[4:0] ? io_in_3_Im : _GEN_1679; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1681 = 5'h4 == _T_184[4:0] ? io_in_4_Im : _GEN_1680; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1682 = 5'h5 == _T_184[4:0] ? io_in_5_Im : _GEN_1681; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1683 = 5'h6 == _T_184[4:0] ? io_in_6_Im : _GEN_1682; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1684 = 5'h7 == _T_184[4:0] ? io_in_7_Im : _GEN_1683; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1685 = 5'h8 == _T_184[4:0] ? io_in_8_Im : _GEN_1684; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1686 = 5'h9 == _T_184[4:0] ? io_in_9_Im : _GEN_1685; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1687 = 5'ha == _T_184[4:0] ? io_in_10_Im : _GEN_1686; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1688 = 5'hb == _T_184[4:0] ? io_in_11_Im : _GEN_1687; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1689 = 5'hc == _T_184[4:0] ? io_in_12_Im : _GEN_1688; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1690 = 5'hd == _T_184[4:0] ? io_in_13_Im : _GEN_1689; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1691 = 5'he == _T_184[4:0] ? io_in_14_Im : _GEN_1690; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1692 = 5'hf == _T_184[4:0] ? io_in_15_Im : _GEN_1691; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1693 = 5'h10 == _T_184[4:0] ? io_in_16_Im : _GEN_1692; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1694 = 5'h11 == _T_184[4:0] ? io_in_17_Im : _GEN_1693; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1695 = 5'h12 == _T_184[4:0] ? io_in_18_Im : _GEN_1694; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1696 = 5'h13 == _T_184[4:0] ? io_in_19_Im : _GEN_1695; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1697 = 5'h14 == _T_184[4:0] ? io_in_20_Im : _GEN_1696; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1698 = 5'h15 == _T_184[4:0] ? io_in_21_Im : _GEN_1697; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1699 = 5'h16 == _T_184[4:0] ? io_in_22_Im : _GEN_1698; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1700 = 5'h17 == _T_184[4:0] ? io_in_23_Im : _GEN_1699; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1701 = 5'h18 == _T_184[4:0] ? io_in_24_Im : _GEN_1700; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1702 = 5'h19 == _T_184[4:0] ? io_in_25_Im : _GEN_1701; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1705 = 5'h1 == _T_184[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1706 = 5'h2 == _T_184[4:0] ? io_in_2_Re : _GEN_1705; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1707 = 5'h3 == _T_184[4:0] ? io_in_3_Re : _GEN_1706; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1708 = 5'h4 == _T_184[4:0] ? io_in_4_Re : _GEN_1707; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1709 = 5'h5 == _T_184[4:0] ? io_in_5_Re : _GEN_1708; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1710 = 5'h6 == _T_184[4:0] ? io_in_6_Re : _GEN_1709; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1711 = 5'h7 == _T_184[4:0] ? io_in_7_Re : _GEN_1710; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1712 = 5'h8 == _T_184[4:0] ? io_in_8_Re : _GEN_1711; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1713 = 5'h9 == _T_184[4:0] ? io_in_9_Re : _GEN_1712; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1714 = 5'ha == _T_184[4:0] ? io_in_10_Re : _GEN_1713; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1715 = 5'hb == _T_184[4:0] ? io_in_11_Re : _GEN_1714; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1716 = 5'hc == _T_184[4:0] ? io_in_12_Re : _GEN_1715; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1717 = 5'hd == _T_184[4:0] ? io_in_13_Re : _GEN_1716; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1718 = 5'he == _T_184[4:0] ? io_in_14_Re : _GEN_1717; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1719 = 5'hf == _T_184[4:0] ? io_in_15_Re : _GEN_1718; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1720 = 5'h10 == _T_184[4:0] ? io_in_16_Re : _GEN_1719; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1721 = 5'h11 == _T_184[4:0] ? io_in_17_Re : _GEN_1720; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1722 = 5'h12 == _T_184[4:0] ? io_in_18_Re : _GEN_1721; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1723 = 5'h13 == _T_184[4:0] ? io_in_19_Re : _GEN_1722; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1724 = 5'h14 == _T_184[4:0] ? io_in_20_Re : _GEN_1723; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1725 = 5'h15 == _T_184[4:0] ? io_in_21_Re : _GEN_1724; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1726 = 5'h16 == _T_184[4:0] ? io_in_22_Re : _GEN_1725; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1727 = 5'h17 == _T_184[4:0] ? io_in_23_Re : _GEN_1726; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1728 = 5'h18 == _T_184[4:0] ? io_in_24_Re : _GEN_1727; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1729 = 5'h19 == _T_184[4:0] ? io_in_25_Re : _GEN_1728; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_196 = _T_2 + 37'h10; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1741 = 5'ha == _T_196[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1742 = 5'hb == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1741; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1743 = 5'hc == _T_196[4:0] ? 32'h3f800000 : _GEN_1742; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1744 = 5'hd == _T_196[4:0] ? 32'h3f441b7c : _GEN_1743; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1745 = 5'he == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1744; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1746 = 5'hf == _T_196[4:0] ? 32'h3f800000 : _GEN_1745; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1747 = 5'h10 == _T_196[4:0] ? 32'h3f441b7c : _GEN_1746; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1748 = 5'h11 == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1747; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1749 = 5'h12 == _T_196[4:0] ? 32'h3f800000 : _GEN_1748; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1750 = 5'h13 == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1749; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1751 = 5'h14 == _T_196[4:0] ? 32'hbf708fb2 : _GEN_1750; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1752 = 5'h15 == _T_196[4:0] ? 32'h3f800000 : _GEN_1751; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1753 = 5'h16 == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1752; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1754 = 5'h17 == _T_196[4:0] ? 32'hbf708fb2 : _GEN_1753; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1755 = 5'h18 == _T_196[4:0] ? 32'h3f800000 : _GEN_1754; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1756 = 5'h19 == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1755; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1768 = 5'ha == _T_196[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1769 = 5'hb == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1768; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1770 = 5'hc == _T_196[4:0] ? 32'h80800000 : _GEN_1769; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1771 = 5'hd == _T_196[4:0] ? 32'hbf248dba : _GEN_1770; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1772 = 5'he == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1771; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1773 = 5'hf == _T_196[4:0] ? 32'h80800000 : _GEN_1772; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1774 = 5'h10 == _T_196[4:0] ? 32'hbf248dba : _GEN_1773; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1775 = 5'h11 == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1774; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1776 = 5'h12 == _T_196[4:0] ? 32'h80800000 : _GEN_1775; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1777 = 5'h13 == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1776; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1778 = 5'h14 == _T_196[4:0] ? 32'hbeaf1d40 : _GEN_1777; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1779 = 5'h15 == _T_196[4:0] ? 32'h80800000 : _GEN_1778; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1780 = 5'h16 == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1779; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1781 = 5'h17 == _T_196[4:0] ? 32'hbeaf1d40 : _GEN_1780; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1782 = 5'h18 == _T_196[4:0] ? 32'h80800000 : _GEN_1781; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1783 = 5'h19 == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1782; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1786 = 5'h1 == _T_196[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1787 = 5'h2 == _T_196[4:0] ? io_in_2_Im : _GEN_1786; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1788 = 5'h3 == _T_196[4:0] ? io_in_3_Im : _GEN_1787; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1789 = 5'h4 == _T_196[4:0] ? io_in_4_Im : _GEN_1788; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1790 = 5'h5 == _T_196[4:0] ? io_in_5_Im : _GEN_1789; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1791 = 5'h6 == _T_196[4:0] ? io_in_6_Im : _GEN_1790; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1792 = 5'h7 == _T_196[4:0] ? io_in_7_Im : _GEN_1791; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1793 = 5'h8 == _T_196[4:0] ? io_in_8_Im : _GEN_1792; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1794 = 5'h9 == _T_196[4:0] ? io_in_9_Im : _GEN_1793; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1795 = 5'ha == _T_196[4:0] ? io_in_10_Im : _GEN_1794; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1796 = 5'hb == _T_196[4:0] ? io_in_11_Im : _GEN_1795; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1797 = 5'hc == _T_196[4:0] ? io_in_12_Im : _GEN_1796; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1798 = 5'hd == _T_196[4:0] ? io_in_13_Im : _GEN_1797; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1799 = 5'he == _T_196[4:0] ? io_in_14_Im : _GEN_1798; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1800 = 5'hf == _T_196[4:0] ? io_in_15_Im : _GEN_1799; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1801 = 5'h10 == _T_196[4:0] ? io_in_16_Im : _GEN_1800; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1802 = 5'h11 == _T_196[4:0] ? io_in_17_Im : _GEN_1801; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1803 = 5'h12 == _T_196[4:0] ? io_in_18_Im : _GEN_1802; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1804 = 5'h13 == _T_196[4:0] ? io_in_19_Im : _GEN_1803; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1805 = 5'h14 == _T_196[4:0] ? io_in_20_Im : _GEN_1804; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1806 = 5'h15 == _T_196[4:0] ? io_in_21_Im : _GEN_1805; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1807 = 5'h16 == _T_196[4:0] ? io_in_22_Im : _GEN_1806; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1808 = 5'h17 == _T_196[4:0] ? io_in_23_Im : _GEN_1807; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1809 = 5'h18 == _T_196[4:0] ? io_in_24_Im : _GEN_1808; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1810 = 5'h19 == _T_196[4:0] ? io_in_25_Im : _GEN_1809; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1813 = 5'h1 == _T_196[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1814 = 5'h2 == _T_196[4:0] ? io_in_2_Re : _GEN_1813; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1815 = 5'h3 == _T_196[4:0] ? io_in_3_Re : _GEN_1814; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1816 = 5'h4 == _T_196[4:0] ? io_in_4_Re : _GEN_1815; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1817 = 5'h5 == _T_196[4:0] ? io_in_5_Re : _GEN_1816; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1818 = 5'h6 == _T_196[4:0] ? io_in_6_Re : _GEN_1817; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1819 = 5'h7 == _T_196[4:0] ? io_in_7_Re : _GEN_1818; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1820 = 5'h8 == _T_196[4:0] ? io_in_8_Re : _GEN_1819; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1821 = 5'h9 == _T_196[4:0] ? io_in_9_Re : _GEN_1820; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1822 = 5'ha == _T_196[4:0] ? io_in_10_Re : _GEN_1821; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1823 = 5'hb == _T_196[4:0] ? io_in_11_Re : _GEN_1822; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1824 = 5'hc == _T_196[4:0] ? io_in_12_Re : _GEN_1823; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1825 = 5'hd == _T_196[4:0] ? io_in_13_Re : _GEN_1824; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1826 = 5'he == _T_196[4:0] ? io_in_14_Re : _GEN_1825; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1827 = 5'hf == _T_196[4:0] ? io_in_15_Re : _GEN_1826; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1828 = 5'h10 == _T_196[4:0] ? io_in_16_Re : _GEN_1827; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1829 = 5'h11 == _T_196[4:0] ? io_in_17_Re : _GEN_1828; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1830 = 5'h12 == _T_196[4:0] ? io_in_18_Re : _GEN_1829; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1831 = 5'h13 == _T_196[4:0] ? io_in_19_Re : _GEN_1830; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1832 = 5'h14 == _T_196[4:0] ? io_in_20_Re : _GEN_1831; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1833 = 5'h15 == _T_196[4:0] ? io_in_21_Re : _GEN_1832; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1834 = 5'h16 == _T_196[4:0] ? io_in_22_Re : _GEN_1833; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1835 = 5'h17 == _T_196[4:0] ? io_in_23_Re : _GEN_1834; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1836 = 5'h18 == _T_196[4:0] ? io_in_24_Re : _GEN_1835; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1837 = 5'h19 == _T_196[4:0] ? io_in_25_Re : _GEN_1836; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_208 = _T_2 + 37'h11; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1849 = 5'ha == _T_208[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1850 = 5'hb == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1849; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1851 = 5'hc == _T_208[4:0] ? 32'h3f800000 : _GEN_1850; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1852 = 5'hd == _T_208[4:0] ? 32'h3f441b7c : _GEN_1851; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1853 = 5'he == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1852; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1854 = 5'hf == _T_208[4:0] ? 32'h3f800000 : _GEN_1853; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1855 = 5'h10 == _T_208[4:0] ? 32'h3f441b7c : _GEN_1854; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1856 = 5'h11 == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1855; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1857 = 5'h12 == _T_208[4:0] ? 32'h3f800000 : _GEN_1856; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1858 = 5'h13 == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1857; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1859 = 5'h14 == _T_208[4:0] ? 32'hbf708fb2 : _GEN_1858; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1860 = 5'h15 == _T_208[4:0] ? 32'h3f800000 : _GEN_1859; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1861 = 5'h16 == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1860; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1862 = 5'h17 == _T_208[4:0] ? 32'hbf708fb2 : _GEN_1861; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1863 = 5'h18 == _T_208[4:0] ? 32'h3f800000 : _GEN_1862; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1864 = 5'h19 == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1863; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1876 = 5'ha == _T_208[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1877 = 5'hb == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1876; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1878 = 5'hc == _T_208[4:0] ? 32'h80800000 : _GEN_1877; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1879 = 5'hd == _T_208[4:0] ? 32'hbf248dba : _GEN_1878; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1880 = 5'he == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1879; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1881 = 5'hf == _T_208[4:0] ? 32'h80800000 : _GEN_1880; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1882 = 5'h10 == _T_208[4:0] ? 32'hbf248dba : _GEN_1881; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1883 = 5'h11 == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1882; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1884 = 5'h12 == _T_208[4:0] ? 32'h80800000 : _GEN_1883; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1885 = 5'h13 == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1884; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1886 = 5'h14 == _T_208[4:0] ? 32'hbeaf1d40 : _GEN_1885; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1887 = 5'h15 == _T_208[4:0] ? 32'h80800000 : _GEN_1886; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1888 = 5'h16 == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1887; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1889 = 5'h17 == _T_208[4:0] ? 32'hbeaf1d40 : _GEN_1888; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1890 = 5'h18 == _T_208[4:0] ? 32'h80800000 : _GEN_1889; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1891 = 5'h19 == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1890; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1894 = 5'h1 == _T_208[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1895 = 5'h2 == _T_208[4:0] ? io_in_2_Im : _GEN_1894; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1896 = 5'h3 == _T_208[4:0] ? io_in_3_Im : _GEN_1895; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1897 = 5'h4 == _T_208[4:0] ? io_in_4_Im : _GEN_1896; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1898 = 5'h5 == _T_208[4:0] ? io_in_5_Im : _GEN_1897; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1899 = 5'h6 == _T_208[4:0] ? io_in_6_Im : _GEN_1898; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1900 = 5'h7 == _T_208[4:0] ? io_in_7_Im : _GEN_1899; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1901 = 5'h8 == _T_208[4:0] ? io_in_8_Im : _GEN_1900; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1902 = 5'h9 == _T_208[4:0] ? io_in_9_Im : _GEN_1901; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1903 = 5'ha == _T_208[4:0] ? io_in_10_Im : _GEN_1902; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1904 = 5'hb == _T_208[4:0] ? io_in_11_Im : _GEN_1903; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1905 = 5'hc == _T_208[4:0] ? io_in_12_Im : _GEN_1904; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1906 = 5'hd == _T_208[4:0] ? io_in_13_Im : _GEN_1905; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1907 = 5'he == _T_208[4:0] ? io_in_14_Im : _GEN_1906; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1908 = 5'hf == _T_208[4:0] ? io_in_15_Im : _GEN_1907; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1909 = 5'h10 == _T_208[4:0] ? io_in_16_Im : _GEN_1908; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1910 = 5'h11 == _T_208[4:0] ? io_in_17_Im : _GEN_1909; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1911 = 5'h12 == _T_208[4:0] ? io_in_18_Im : _GEN_1910; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1912 = 5'h13 == _T_208[4:0] ? io_in_19_Im : _GEN_1911; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1913 = 5'h14 == _T_208[4:0] ? io_in_20_Im : _GEN_1912; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1914 = 5'h15 == _T_208[4:0] ? io_in_21_Im : _GEN_1913; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1915 = 5'h16 == _T_208[4:0] ? io_in_22_Im : _GEN_1914; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1916 = 5'h17 == _T_208[4:0] ? io_in_23_Im : _GEN_1915; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1917 = 5'h18 == _T_208[4:0] ? io_in_24_Im : _GEN_1916; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1918 = 5'h19 == _T_208[4:0] ? io_in_25_Im : _GEN_1917; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1921 = 5'h1 == _T_208[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1922 = 5'h2 == _T_208[4:0] ? io_in_2_Re : _GEN_1921; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1923 = 5'h3 == _T_208[4:0] ? io_in_3_Re : _GEN_1922; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1924 = 5'h4 == _T_208[4:0] ? io_in_4_Re : _GEN_1923; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1925 = 5'h5 == _T_208[4:0] ? io_in_5_Re : _GEN_1924; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1926 = 5'h6 == _T_208[4:0] ? io_in_6_Re : _GEN_1925; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1927 = 5'h7 == _T_208[4:0] ? io_in_7_Re : _GEN_1926; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1928 = 5'h8 == _T_208[4:0] ? io_in_8_Re : _GEN_1927; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1929 = 5'h9 == _T_208[4:0] ? io_in_9_Re : _GEN_1928; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1930 = 5'ha == _T_208[4:0] ? io_in_10_Re : _GEN_1929; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1931 = 5'hb == _T_208[4:0] ? io_in_11_Re : _GEN_1930; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1932 = 5'hc == _T_208[4:0] ? io_in_12_Re : _GEN_1931; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1933 = 5'hd == _T_208[4:0] ? io_in_13_Re : _GEN_1932; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1934 = 5'he == _T_208[4:0] ? io_in_14_Re : _GEN_1933; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1935 = 5'hf == _T_208[4:0] ? io_in_15_Re : _GEN_1934; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1936 = 5'h10 == _T_208[4:0] ? io_in_16_Re : _GEN_1935; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1937 = 5'h11 == _T_208[4:0] ? io_in_17_Re : _GEN_1936; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1938 = 5'h12 == _T_208[4:0] ? io_in_18_Re : _GEN_1937; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1939 = 5'h13 == _T_208[4:0] ? io_in_19_Re : _GEN_1938; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1940 = 5'h14 == _T_208[4:0] ? io_in_20_Re : _GEN_1939; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1941 = 5'h15 == _T_208[4:0] ? io_in_21_Re : _GEN_1940; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1942 = 5'h16 == _T_208[4:0] ? io_in_22_Re : _GEN_1941; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1943 = 5'h17 == _T_208[4:0] ? io_in_23_Re : _GEN_1942; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1944 = 5'h18 == _T_208[4:0] ? io_in_24_Re : _GEN_1943; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1945 = 5'h19 == _T_208[4:0] ? io_in_25_Re : _GEN_1944; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_220 = _T_2 + 37'h12; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1957 = 5'ha == _T_220[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1958 = 5'hb == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1957; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1959 = 5'hc == _T_220[4:0] ? 32'h3f800000 : _GEN_1958; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1960 = 5'hd == _T_220[4:0] ? 32'h3f441b7c : _GEN_1959; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1961 = 5'he == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1960; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1962 = 5'hf == _T_220[4:0] ? 32'h3f800000 : _GEN_1961; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1963 = 5'h10 == _T_220[4:0] ? 32'h3f441b7c : _GEN_1962; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1964 = 5'h11 == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1963; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1965 = 5'h12 == _T_220[4:0] ? 32'h3f800000 : _GEN_1964; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1966 = 5'h13 == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1965; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1967 = 5'h14 == _T_220[4:0] ? 32'hbf708fb2 : _GEN_1966; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1968 = 5'h15 == _T_220[4:0] ? 32'h3f800000 : _GEN_1967; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1969 = 5'h16 == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1968; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1970 = 5'h17 == _T_220[4:0] ? 32'hbf708fb2 : _GEN_1969; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1971 = 5'h18 == _T_220[4:0] ? 32'h3f800000 : _GEN_1970; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1972 = 5'h19 == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1971; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1984 = 5'ha == _T_220[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1985 = 5'hb == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1984; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1986 = 5'hc == _T_220[4:0] ? 32'h80800000 : _GEN_1985; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1987 = 5'hd == _T_220[4:0] ? 32'hbf248dba : _GEN_1986; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1988 = 5'he == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1987; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1989 = 5'hf == _T_220[4:0] ? 32'h80800000 : _GEN_1988; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1990 = 5'h10 == _T_220[4:0] ? 32'hbf248dba : _GEN_1989; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1991 = 5'h11 == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1990; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1992 = 5'h12 == _T_220[4:0] ? 32'h80800000 : _GEN_1991; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1993 = 5'h13 == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1992; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1994 = 5'h14 == _T_220[4:0] ? 32'hbeaf1d40 : _GEN_1993; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1995 = 5'h15 == _T_220[4:0] ? 32'h80800000 : _GEN_1994; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1996 = 5'h16 == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1995; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1997 = 5'h17 == _T_220[4:0] ? 32'hbeaf1d40 : _GEN_1996; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1998 = 5'h18 == _T_220[4:0] ? 32'h80800000 : _GEN_1997; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1999 = 5'h19 == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1998; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2002 = 5'h1 == _T_220[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2003 = 5'h2 == _T_220[4:0] ? io_in_2_Im : _GEN_2002; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2004 = 5'h3 == _T_220[4:0] ? io_in_3_Im : _GEN_2003; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2005 = 5'h4 == _T_220[4:0] ? io_in_4_Im : _GEN_2004; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2006 = 5'h5 == _T_220[4:0] ? io_in_5_Im : _GEN_2005; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2007 = 5'h6 == _T_220[4:0] ? io_in_6_Im : _GEN_2006; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2008 = 5'h7 == _T_220[4:0] ? io_in_7_Im : _GEN_2007; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2009 = 5'h8 == _T_220[4:0] ? io_in_8_Im : _GEN_2008; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2010 = 5'h9 == _T_220[4:0] ? io_in_9_Im : _GEN_2009; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2011 = 5'ha == _T_220[4:0] ? io_in_10_Im : _GEN_2010; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2012 = 5'hb == _T_220[4:0] ? io_in_11_Im : _GEN_2011; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2013 = 5'hc == _T_220[4:0] ? io_in_12_Im : _GEN_2012; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2014 = 5'hd == _T_220[4:0] ? io_in_13_Im : _GEN_2013; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2015 = 5'he == _T_220[4:0] ? io_in_14_Im : _GEN_2014; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2016 = 5'hf == _T_220[4:0] ? io_in_15_Im : _GEN_2015; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2017 = 5'h10 == _T_220[4:0] ? io_in_16_Im : _GEN_2016; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2018 = 5'h11 == _T_220[4:0] ? io_in_17_Im : _GEN_2017; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2019 = 5'h12 == _T_220[4:0] ? io_in_18_Im : _GEN_2018; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2020 = 5'h13 == _T_220[4:0] ? io_in_19_Im : _GEN_2019; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2021 = 5'h14 == _T_220[4:0] ? io_in_20_Im : _GEN_2020; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2022 = 5'h15 == _T_220[4:0] ? io_in_21_Im : _GEN_2021; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2023 = 5'h16 == _T_220[4:0] ? io_in_22_Im : _GEN_2022; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2024 = 5'h17 == _T_220[4:0] ? io_in_23_Im : _GEN_2023; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2025 = 5'h18 == _T_220[4:0] ? io_in_24_Im : _GEN_2024; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2026 = 5'h19 == _T_220[4:0] ? io_in_25_Im : _GEN_2025; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2029 = 5'h1 == _T_220[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2030 = 5'h2 == _T_220[4:0] ? io_in_2_Re : _GEN_2029; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2031 = 5'h3 == _T_220[4:0] ? io_in_3_Re : _GEN_2030; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2032 = 5'h4 == _T_220[4:0] ? io_in_4_Re : _GEN_2031; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2033 = 5'h5 == _T_220[4:0] ? io_in_5_Re : _GEN_2032; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2034 = 5'h6 == _T_220[4:0] ? io_in_6_Re : _GEN_2033; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2035 = 5'h7 == _T_220[4:0] ? io_in_7_Re : _GEN_2034; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2036 = 5'h8 == _T_220[4:0] ? io_in_8_Re : _GEN_2035; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2037 = 5'h9 == _T_220[4:0] ? io_in_9_Re : _GEN_2036; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2038 = 5'ha == _T_220[4:0] ? io_in_10_Re : _GEN_2037; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2039 = 5'hb == _T_220[4:0] ? io_in_11_Re : _GEN_2038; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2040 = 5'hc == _T_220[4:0] ? io_in_12_Re : _GEN_2039; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2041 = 5'hd == _T_220[4:0] ? io_in_13_Re : _GEN_2040; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2042 = 5'he == _T_220[4:0] ? io_in_14_Re : _GEN_2041; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2043 = 5'hf == _T_220[4:0] ? io_in_15_Re : _GEN_2042; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2044 = 5'h10 == _T_220[4:0] ? io_in_16_Re : _GEN_2043; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2045 = 5'h11 == _T_220[4:0] ? io_in_17_Re : _GEN_2044; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2046 = 5'h12 == _T_220[4:0] ? io_in_18_Re : _GEN_2045; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2047 = 5'h13 == _T_220[4:0] ? io_in_19_Re : _GEN_2046; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2048 = 5'h14 == _T_220[4:0] ? io_in_20_Re : _GEN_2047; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2049 = 5'h15 == _T_220[4:0] ? io_in_21_Re : _GEN_2048; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2050 = 5'h16 == _T_220[4:0] ? io_in_22_Re : _GEN_2049; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2051 = 5'h17 == _T_220[4:0] ? io_in_23_Re : _GEN_2050; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2052 = 5'h18 == _T_220[4:0] ? io_in_24_Re : _GEN_2051; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2053 = 5'h19 == _T_220[4:0] ? io_in_25_Re : _GEN_2052; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_232 = _T_2 + 37'h13; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2065 = 5'ha == _T_232[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2066 = 5'hb == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2065; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2067 = 5'hc == _T_232[4:0] ? 32'h3f800000 : _GEN_2066; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2068 = 5'hd == _T_232[4:0] ? 32'h3f441b7c : _GEN_2067; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2069 = 5'he == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2068; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2070 = 5'hf == _T_232[4:0] ? 32'h3f800000 : _GEN_2069; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2071 = 5'h10 == _T_232[4:0] ? 32'h3f441b7c : _GEN_2070; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2072 = 5'h11 == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2071; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2073 = 5'h12 == _T_232[4:0] ? 32'h3f800000 : _GEN_2072; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2074 = 5'h13 == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2073; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2075 = 5'h14 == _T_232[4:0] ? 32'hbf708fb2 : _GEN_2074; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2076 = 5'h15 == _T_232[4:0] ? 32'h3f800000 : _GEN_2075; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2077 = 5'h16 == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2076; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2078 = 5'h17 == _T_232[4:0] ? 32'hbf708fb2 : _GEN_2077; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2079 = 5'h18 == _T_232[4:0] ? 32'h3f800000 : _GEN_2078; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2080 = 5'h19 == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2079; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2092 = 5'ha == _T_232[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2093 = 5'hb == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2092; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2094 = 5'hc == _T_232[4:0] ? 32'h80800000 : _GEN_2093; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2095 = 5'hd == _T_232[4:0] ? 32'hbf248dba : _GEN_2094; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2096 = 5'he == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2095; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2097 = 5'hf == _T_232[4:0] ? 32'h80800000 : _GEN_2096; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2098 = 5'h10 == _T_232[4:0] ? 32'hbf248dba : _GEN_2097; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2099 = 5'h11 == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2098; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2100 = 5'h12 == _T_232[4:0] ? 32'h80800000 : _GEN_2099; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2101 = 5'h13 == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2100; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2102 = 5'h14 == _T_232[4:0] ? 32'hbeaf1d40 : _GEN_2101; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2103 = 5'h15 == _T_232[4:0] ? 32'h80800000 : _GEN_2102; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2104 = 5'h16 == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2103; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2105 = 5'h17 == _T_232[4:0] ? 32'hbeaf1d40 : _GEN_2104; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2106 = 5'h18 == _T_232[4:0] ? 32'h80800000 : _GEN_2105; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2107 = 5'h19 == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2106; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2110 = 5'h1 == _T_232[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2111 = 5'h2 == _T_232[4:0] ? io_in_2_Im : _GEN_2110; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2112 = 5'h3 == _T_232[4:0] ? io_in_3_Im : _GEN_2111; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2113 = 5'h4 == _T_232[4:0] ? io_in_4_Im : _GEN_2112; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2114 = 5'h5 == _T_232[4:0] ? io_in_5_Im : _GEN_2113; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2115 = 5'h6 == _T_232[4:0] ? io_in_6_Im : _GEN_2114; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2116 = 5'h7 == _T_232[4:0] ? io_in_7_Im : _GEN_2115; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2117 = 5'h8 == _T_232[4:0] ? io_in_8_Im : _GEN_2116; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2118 = 5'h9 == _T_232[4:0] ? io_in_9_Im : _GEN_2117; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2119 = 5'ha == _T_232[4:0] ? io_in_10_Im : _GEN_2118; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2120 = 5'hb == _T_232[4:0] ? io_in_11_Im : _GEN_2119; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2121 = 5'hc == _T_232[4:0] ? io_in_12_Im : _GEN_2120; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2122 = 5'hd == _T_232[4:0] ? io_in_13_Im : _GEN_2121; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2123 = 5'he == _T_232[4:0] ? io_in_14_Im : _GEN_2122; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2124 = 5'hf == _T_232[4:0] ? io_in_15_Im : _GEN_2123; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2125 = 5'h10 == _T_232[4:0] ? io_in_16_Im : _GEN_2124; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2126 = 5'h11 == _T_232[4:0] ? io_in_17_Im : _GEN_2125; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2127 = 5'h12 == _T_232[4:0] ? io_in_18_Im : _GEN_2126; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2128 = 5'h13 == _T_232[4:0] ? io_in_19_Im : _GEN_2127; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2129 = 5'h14 == _T_232[4:0] ? io_in_20_Im : _GEN_2128; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2130 = 5'h15 == _T_232[4:0] ? io_in_21_Im : _GEN_2129; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2131 = 5'h16 == _T_232[4:0] ? io_in_22_Im : _GEN_2130; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2132 = 5'h17 == _T_232[4:0] ? io_in_23_Im : _GEN_2131; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2133 = 5'h18 == _T_232[4:0] ? io_in_24_Im : _GEN_2132; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2134 = 5'h19 == _T_232[4:0] ? io_in_25_Im : _GEN_2133; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2137 = 5'h1 == _T_232[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2138 = 5'h2 == _T_232[4:0] ? io_in_2_Re : _GEN_2137; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2139 = 5'h3 == _T_232[4:0] ? io_in_3_Re : _GEN_2138; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2140 = 5'h4 == _T_232[4:0] ? io_in_4_Re : _GEN_2139; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2141 = 5'h5 == _T_232[4:0] ? io_in_5_Re : _GEN_2140; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2142 = 5'h6 == _T_232[4:0] ? io_in_6_Re : _GEN_2141; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2143 = 5'h7 == _T_232[4:0] ? io_in_7_Re : _GEN_2142; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2144 = 5'h8 == _T_232[4:0] ? io_in_8_Re : _GEN_2143; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2145 = 5'h9 == _T_232[4:0] ? io_in_9_Re : _GEN_2144; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2146 = 5'ha == _T_232[4:0] ? io_in_10_Re : _GEN_2145; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2147 = 5'hb == _T_232[4:0] ? io_in_11_Re : _GEN_2146; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2148 = 5'hc == _T_232[4:0] ? io_in_12_Re : _GEN_2147; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2149 = 5'hd == _T_232[4:0] ? io_in_13_Re : _GEN_2148; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2150 = 5'he == _T_232[4:0] ? io_in_14_Re : _GEN_2149; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2151 = 5'hf == _T_232[4:0] ? io_in_15_Re : _GEN_2150; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2152 = 5'h10 == _T_232[4:0] ? io_in_16_Re : _GEN_2151; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2153 = 5'h11 == _T_232[4:0] ? io_in_17_Re : _GEN_2152; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2154 = 5'h12 == _T_232[4:0] ? io_in_18_Re : _GEN_2153; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2155 = 5'h13 == _T_232[4:0] ? io_in_19_Re : _GEN_2154; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2156 = 5'h14 == _T_232[4:0] ? io_in_20_Re : _GEN_2155; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2157 = 5'h15 == _T_232[4:0] ? io_in_21_Re : _GEN_2156; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2158 = 5'h16 == _T_232[4:0] ? io_in_22_Re : _GEN_2157; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2159 = 5'h17 == _T_232[4:0] ? io_in_23_Re : _GEN_2158; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2160 = 5'h18 == _T_232[4:0] ? io_in_24_Re : _GEN_2159; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2161 = 5'h19 == _T_232[4:0] ? io_in_25_Re : _GEN_2160; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_244 = _T_2 + 37'h14; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2173 = 5'ha == _T_244[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2174 = 5'hb == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2173; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2175 = 5'hc == _T_244[4:0] ? 32'h3f800000 : _GEN_2174; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2176 = 5'hd == _T_244[4:0] ? 32'h3f441b7c : _GEN_2175; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2177 = 5'he == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2176; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2178 = 5'hf == _T_244[4:0] ? 32'h3f800000 : _GEN_2177; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2179 = 5'h10 == _T_244[4:0] ? 32'h3f441b7c : _GEN_2178; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2180 = 5'h11 == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2179; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2181 = 5'h12 == _T_244[4:0] ? 32'h3f800000 : _GEN_2180; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2182 = 5'h13 == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2181; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2183 = 5'h14 == _T_244[4:0] ? 32'hbf708fb2 : _GEN_2182; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2184 = 5'h15 == _T_244[4:0] ? 32'h3f800000 : _GEN_2183; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2185 = 5'h16 == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2184; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2186 = 5'h17 == _T_244[4:0] ? 32'hbf708fb2 : _GEN_2185; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2187 = 5'h18 == _T_244[4:0] ? 32'h3f800000 : _GEN_2186; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2188 = 5'h19 == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2187; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2200 = 5'ha == _T_244[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2201 = 5'hb == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2200; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2202 = 5'hc == _T_244[4:0] ? 32'h80800000 : _GEN_2201; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2203 = 5'hd == _T_244[4:0] ? 32'hbf248dba : _GEN_2202; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2204 = 5'he == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2203; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2205 = 5'hf == _T_244[4:0] ? 32'h80800000 : _GEN_2204; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2206 = 5'h10 == _T_244[4:0] ? 32'hbf248dba : _GEN_2205; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2207 = 5'h11 == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2206; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2208 = 5'h12 == _T_244[4:0] ? 32'h80800000 : _GEN_2207; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2209 = 5'h13 == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2208; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2210 = 5'h14 == _T_244[4:0] ? 32'hbeaf1d40 : _GEN_2209; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2211 = 5'h15 == _T_244[4:0] ? 32'h80800000 : _GEN_2210; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2212 = 5'h16 == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2211; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2213 = 5'h17 == _T_244[4:0] ? 32'hbeaf1d40 : _GEN_2212; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2214 = 5'h18 == _T_244[4:0] ? 32'h80800000 : _GEN_2213; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2215 = 5'h19 == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2214; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2218 = 5'h1 == _T_244[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2219 = 5'h2 == _T_244[4:0] ? io_in_2_Im : _GEN_2218; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2220 = 5'h3 == _T_244[4:0] ? io_in_3_Im : _GEN_2219; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2221 = 5'h4 == _T_244[4:0] ? io_in_4_Im : _GEN_2220; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2222 = 5'h5 == _T_244[4:0] ? io_in_5_Im : _GEN_2221; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2223 = 5'h6 == _T_244[4:0] ? io_in_6_Im : _GEN_2222; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2224 = 5'h7 == _T_244[4:0] ? io_in_7_Im : _GEN_2223; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2225 = 5'h8 == _T_244[4:0] ? io_in_8_Im : _GEN_2224; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2226 = 5'h9 == _T_244[4:0] ? io_in_9_Im : _GEN_2225; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2227 = 5'ha == _T_244[4:0] ? io_in_10_Im : _GEN_2226; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2228 = 5'hb == _T_244[4:0] ? io_in_11_Im : _GEN_2227; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2229 = 5'hc == _T_244[4:0] ? io_in_12_Im : _GEN_2228; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2230 = 5'hd == _T_244[4:0] ? io_in_13_Im : _GEN_2229; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2231 = 5'he == _T_244[4:0] ? io_in_14_Im : _GEN_2230; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2232 = 5'hf == _T_244[4:0] ? io_in_15_Im : _GEN_2231; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2233 = 5'h10 == _T_244[4:0] ? io_in_16_Im : _GEN_2232; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2234 = 5'h11 == _T_244[4:0] ? io_in_17_Im : _GEN_2233; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2235 = 5'h12 == _T_244[4:0] ? io_in_18_Im : _GEN_2234; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2236 = 5'h13 == _T_244[4:0] ? io_in_19_Im : _GEN_2235; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2237 = 5'h14 == _T_244[4:0] ? io_in_20_Im : _GEN_2236; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2238 = 5'h15 == _T_244[4:0] ? io_in_21_Im : _GEN_2237; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2239 = 5'h16 == _T_244[4:0] ? io_in_22_Im : _GEN_2238; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2240 = 5'h17 == _T_244[4:0] ? io_in_23_Im : _GEN_2239; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2241 = 5'h18 == _T_244[4:0] ? io_in_24_Im : _GEN_2240; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2242 = 5'h19 == _T_244[4:0] ? io_in_25_Im : _GEN_2241; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2245 = 5'h1 == _T_244[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2246 = 5'h2 == _T_244[4:0] ? io_in_2_Re : _GEN_2245; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2247 = 5'h3 == _T_244[4:0] ? io_in_3_Re : _GEN_2246; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2248 = 5'h4 == _T_244[4:0] ? io_in_4_Re : _GEN_2247; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2249 = 5'h5 == _T_244[4:0] ? io_in_5_Re : _GEN_2248; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2250 = 5'h6 == _T_244[4:0] ? io_in_6_Re : _GEN_2249; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2251 = 5'h7 == _T_244[4:0] ? io_in_7_Re : _GEN_2250; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2252 = 5'h8 == _T_244[4:0] ? io_in_8_Re : _GEN_2251; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2253 = 5'h9 == _T_244[4:0] ? io_in_9_Re : _GEN_2252; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2254 = 5'ha == _T_244[4:0] ? io_in_10_Re : _GEN_2253; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2255 = 5'hb == _T_244[4:0] ? io_in_11_Re : _GEN_2254; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2256 = 5'hc == _T_244[4:0] ? io_in_12_Re : _GEN_2255; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2257 = 5'hd == _T_244[4:0] ? io_in_13_Re : _GEN_2256; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2258 = 5'he == _T_244[4:0] ? io_in_14_Re : _GEN_2257; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2259 = 5'hf == _T_244[4:0] ? io_in_15_Re : _GEN_2258; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2260 = 5'h10 == _T_244[4:0] ? io_in_16_Re : _GEN_2259; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2261 = 5'h11 == _T_244[4:0] ? io_in_17_Re : _GEN_2260; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2262 = 5'h12 == _T_244[4:0] ? io_in_18_Re : _GEN_2261; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2263 = 5'h13 == _T_244[4:0] ? io_in_19_Re : _GEN_2262; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2264 = 5'h14 == _T_244[4:0] ? io_in_20_Re : _GEN_2263; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2265 = 5'h15 == _T_244[4:0] ? io_in_21_Re : _GEN_2264; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2266 = 5'h16 == _T_244[4:0] ? io_in_22_Re : _GEN_2265; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2267 = 5'h17 == _T_244[4:0] ? io_in_23_Re : _GEN_2266; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2268 = 5'h18 == _T_244[4:0] ? io_in_24_Re : _GEN_2267; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2269 = 5'h19 == _T_244[4:0] ? io_in_25_Re : _GEN_2268; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_256 = _T_2 + 37'h15; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2281 = 5'ha == _T_256[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2282 = 5'hb == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2281; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2283 = 5'hc == _T_256[4:0] ? 32'h3f800000 : _GEN_2282; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2284 = 5'hd == _T_256[4:0] ? 32'h3f441b7c : _GEN_2283; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2285 = 5'he == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2284; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2286 = 5'hf == _T_256[4:0] ? 32'h3f800000 : _GEN_2285; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2287 = 5'h10 == _T_256[4:0] ? 32'h3f441b7c : _GEN_2286; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2288 = 5'h11 == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2287; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2289 = 5'h12 == _T_256[4:0] ? 32'h3f800000 : _GEN_2288; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2290 = 5'h13 == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2289; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2291 = 5'h14 == _T_256[4:0] ? 32'hbf708fb2 : _GEN_2290; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2292 = 5'h15 == _T_256[4:0] ? 32'h3f800000 : _GEN_2291; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2293 = 5'h16 == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2292; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2294 = 5'h17 == _T_256[4:0] ? 32'hbf708fb2 : _GEN_2293; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2295 = 5'h18 == _T_256[4:0] ? 32'h3f800000 : _GEN_2294; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2296 = 5'h19 == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2295; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2308 = 5'ha == _T_256[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2309 = 5'hb == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2308; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2310 = 5'hc == _T_256[4:0] ? 32'h80800000 : _GEN_2309; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2311 = 5'hd == _T_256[4:0] ? 32'hbf248dba : _GEN_2310; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2312 = 5'he == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2311; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2313 = 5'hf == _T_256[4:0] ? 32'h80800000 : _GEN_2312; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2314 = 5'h10 == _T_256[4:0] ? 32'hbf248dba : _GEN_2313; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2315 = 5'h11 == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2314; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2316 = 5'h12 == _T_256[4:0] ? 32'h80800000 : _GEN_2315; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2317 = 5'h13 == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2316; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2318 = 5'h14 == _T_256[4:0] ? 32'hbeaf1d40 : _GEN_2317; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2319 = 5'h15 == _T_256[4:0] ? 32'h80800000 : _GEN_2318; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2320 = 5'h16 == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2319; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2321 = 5'h17 == _T_256[4:0] ? 32'hbeaf1d40 : _GEN_2320; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2322 = 5'h18 == _T_256[4:0] ? 32'h80800000 : _GEN_2321; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2323 = 5'h19 == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2322; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2326 = 5'h1 == _T_256[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2327 = 5'h2 == _T_256[4:0] ? io_in_2_Im : _GEN_2326; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2328 = 5'h3 == _T_256[4:0] ? io_in_3_Im : _GEN_2327; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2329 = 5'h4 == _T_256[4:0] ? io_in_4_Im : _GEN_2328; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2330 = 5'h5 == _T_256[4:0] ? io_in_5_Im : _GEN_2329; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2331 = 5'h6 == _T_256[4:0] ? io_in_6_Im : _GEN_2330; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2332 = 5'h7 == _T_256[4:0] ? io_in_7_Im : _GEN_2331; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2333 = 5'h8 == _T_256[4:0] ? io_in_8_Im : _GEN_2332; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2334 = 5'h9 == _T_256[4:0] ? io_in_9_Im : _GEN_2333; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2335 = 5'ha == _T_256[4:0] ? io_in_10_Im : _GEN_2334; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2336 = 5'hb == _T_256[4:0] ? io_in_11_Im : _GEN_2335; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2337 = 5'hc == _T_256[4:0] ? io_in_12_Im : _GEN_2336; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2338 = 5'hd == _T_256[4:0] ? io_in_13_Im : _GEN_2337; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2339 = 5'he == _T_256[4:0] ? io_in_14_Im : _GEN_2338; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2340 = 5'hf == _T_256[4:0] ? io_in_15_Im : _GEN_2339; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2341 = 5'h10 == _T_256[4:0] ? io_in_16_Im : _GEN_2340; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2342 = 5'h11 == _T_256[4:0] ? io_in_17_Im : _GEN_2341; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2343 = 5'h12 == _T_256[4:0] ? io_in_18_Im : _GEN_2342; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2344 = 5'h13 == _T_256[4:0] ? io_in_19_Im : _GEN_2343; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2345 = 5'h14 == _T_256[4:0] ? io_in_20_Im : _GEN_2344; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2346 = 5'h15 == _T_256[4:0] ? io_in_21_Im : _GEN_2345; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2347 = 5'h16 == _T_256[4:0] ? io_in_22_Im : _GEN_2346; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2348 = 5'h17 == _T_256[4:0] ? io_in_23_Im : _GEN_2347; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2349 = 5'h18 == _T_256[4:0] ? io_in_24_Im : _GEN_2348; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2350 = 5'h19 == _T_256[4:0] ? io_in_25_Im : _GEN_2349; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2353 = 5'h1 == _T_256[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2354 = 5'h2 == _T_256[4:0] ? io_in_2_Re : _GEN_2353; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2355 = 5'h3 == _T_256[4:0] ? io_in_3_Re : _GEN_2354; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2356 = 5'h4 == _T_256[4:0] ? io_in_4_Re : _GEN_2355; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2357 = 5'h5 == _T_256[4:0] ? io_in_5_Re : _GEN_2356; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2358 = 5'h6 == _T_256[4:0] ? io_in_6_Re : _GEN_2357; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2359 = 5'h7 == _T_256[4:0] ? io_in_7_Re : _GEN_2358; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2360 = 5'h8 == _T_256[4:0] ? io_in_8_Re : _GEN_2359; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2361 = 5'h9 == _T_256[4:0] ? io_in_9_Re : _GEN_2360; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2362 = 5'ha == _T_256[4:0] ? io_in_10_Re : _GEN_2361; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2363 = 5'hb == _T_256[4:0] ? io_in_11_Re : _GEN_2362; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2364 = 5'hc == _T_256[4:0] ? io_in_12_Re : _GEN_2363; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2365 = 5'hd == _T_256[4:0] ? io_in_13_Re : _GEN_2364; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2366 = 5'he == _T_256[4:0] ? io_in_14_Re : _GEN_2365; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2367 = 5'hf == _T_256[4:0] ? io_in_15_Re : _GEN_2366; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2368 = 5'h10 == _T_256[4:0] ? io_in_16_Re : _GEN_2367; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2369 = 5'h11 == _T_256[4:0] ? io_in_17_Re : _GEN_2368; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2370 = 5'h12 == _T_256[4:0] ? io_in_18_Re : _GEN_2369; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2371 = 5'h13 == _T_256[4:0] ? io_in_19_Re : _GEN_2370; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2372 = 5'h14 == _T_256[4:0] ? io_in_20_Re : _GEN_2371; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2373 = 5'h15 == _T_256[4:0] ? io_in_21_Re : _GEN_2372; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2374 = 5'h16 == _T_256[4:0] ? io_in_22_Re : _GEN_2373; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2375 = 5'h17 == _T_256[4:0] ? io_in_23_Re : _GEN_2374; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2376 = 5'h18 == _T_256[4:0] ? io_in_24_Re : _GEN_2375; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2377 = 5'h19 == _T_256[4:0] ? io_in_25_Re : _GEN_2376; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_268 = _T_2 + 37'h16; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2389 = 5'ha == _T_268[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2390 = 5'hb == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2389; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2391 = 5'hc == _T_268[4:0] ? 32'h3f800000 : _GEN_2390; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2392 = 5'hd == _T_268[4:0] ? 32'h3f441b7c : _GEN_2391; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2393 = 5'he == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2392; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2394 = 5'hf == _T_268[4:0] ? 32'h3f800000 : _GEN_2393; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2395 = 5'h10 == _T_268[4:0] ? 32'h3f441b7c : _GEN_2394; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2396 = 5'h11 == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2395; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2397 = 5'h12 == _T_268[4:0] ? 32'h3f800000 : _GEN_2396; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2398 = 5'h13 == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2397; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2399 = 5'h14 == _T_268[4:0] ? 32'hbf708fb2 : _GEN_2398; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2400 = 5'h15 == _T_268[4:0] ? 32'h3f800000 : _GEN_2399; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2401 = 5'h16 == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2400; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2402 = 5'h17 == _T_268[4:0] ? 32'hbf708fb2 : _GEN_2401; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2403 = 5'h18 == _T_268[4:0] ? 32'h3f800000 : _GEN_2402; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2404 = 5'h19 == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2403; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2416 = 5'ha == _T_268[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2417 = 5'hb == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2416; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2418 = 5'hc == _T_268[4:0] ? 32'h80800000 : _GEN_2417; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2419 = 5'hd == _T_268[4:0] ? 32'hbf248dba : _GEN_2418; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2420 = 5'he == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2419; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2421 = 5'hf == _T_268[4:0] ? 32'h80800000 : _GEN_2420; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2422 = 5'h10 == _T_268[4:0] ? 32'hbf248dba : _GEN_2421; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2423 = 5'h11 == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2422; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2424 = 5'h12 == _T_268[4:0] ? 32'h80800000 : _GEN_2423; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2425 = 5'h13 == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2424; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2426 = 5'h14 == _T_268[4:0] ? 32'hbeaf1d40 : _GEN_2425; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2427 = 5'h15 == _T_268[4:0] ? 32'h80800000 : _GEN_2426; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2428 = 5'h16 == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2427; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2429 = 5'h17 == _T_268[4:0] ? 32'hbeaf1d40 : _GEN_2428; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2430 = 5'h18 == _T_268[4:0] ? 32'h80800000 : _GEN_2429; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2431 = 5'h19 == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2430; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2434 = 5'h1 == _T_268[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2435 = 5'h2 == _T_268[4:0] ? io_in_2_Im : _GEN_2434; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2436 = 5'h3 == _T_268[4:0] ? io_in_3_Im : _GEN_2435; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2437 = 5'h4 == _T_268[4:0] ? io_in_4_Im : _GEN_2436; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2438 = 5'h5 == _T_268[4:0] ? io_in_5_Im : _GEN_2437; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2439 = 5'h6 == _T_268[4:0] ? io_in_6_Im : _GEN_2438; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2440 = 5'h7 == _T_268[4:0] ? io_in_7_Im : _GEN_2439; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2441 = 5'h8 == _T_268[4:0] ? io_in_8_Im : _GEN_2440; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2442 = 5'h9 == _T_268[4:0] ? io_in_9_Im : _GEN_2441; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2443 = 5'ha == _T_268[4:0] ? io_in_10_Im : _GEN_2442; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2444 = 5'hb == _T_268[4:0] ? io_in_11_Im : _GEN_2443; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2445 = 5'hc == _T_268[4:0] ? io_in_12_Im : _GEN_2444; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2446 = 5'hd == _T_268[4:0] ? io_in_13_Im : _GEN_2445; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2447 = 5'he == _T_268[4:0] ? io_in_14_Im : _GEN_2446; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2448 = 5'hf == _T_268[4:0] ? io_in_15_Im : _GEN_2447; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2449 = 5'h10 == _T_268[4:0] ? io_in_16_Im : _GEN_2448; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2450 = 5'h11 == _T_268[4:0] ? io_in_17_Im : _GEN_2449; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2451 = 5'h12 == _T_268[4:0] ? io_in_18_Im : _GEN_2450; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2452 = 5'h13 == _T_268[4:0] ? io_in_19_Im : _GEN_2451; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2453 = 5'h14 == _T_268[4:0] ? io_in_20_Im : _GEN_2452; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2454 = 5'h15 == _T_268[4:0] ? io_in_21_Im : _GEN_2453; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2455 = 5'h16 == _T_268[4:0] ? io_in_22_Im : _GEN_2454; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2456 = 5'h17 == _T_268[4:0] ? io_in_23_Im : _GEN_2455; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2457 = 5'h18 == _T_268[4:0] ? io_in_24_Im : _GEN_2456; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2458 = 5'h19 == _T_268[4:0] ? io_in_25_Im : _GEN_2457; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2461 = 5'h1 == _T_268[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2462 = 5'h2 == _T_268[4:0] ? io_in_2_Re : _GEN_2461; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2463 = 5'h3 == _T_268[4:0] ? io_in_3_Re : _GEN_2462; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2464 = 5'h4 == _T_268[4:0] ? io_in_4_Re : _GEN_2463; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2465 = 5'h5 == _T_268[4:0] ? io_in_5_Re : _GEN_2464; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2466 = 5'h6 == _T_268[4:0] ? io_in_6_Re : _GEN_2465; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2467 = 5'h7 == _T_268[4:0] ? io_in_7_Re : _GEN_2466; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2468 = 5'h8 == _T_268[4:0] ? io_in_8_Re : _GEN_2467; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2469 = 5'h9 == _T_268[4:0] ? io_in_9_Re : _GEN_2468; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2470 = 5'ha == _T_268[4:0] ? io_in_10_Re : _GEN_2469; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2471 = 5'hb == _T_268[4:0] ? io_in_11_Re : _GEN_2470; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2472 = 5'hc == _T_268[4:0] ? io_in_12_Re : _GEN_2471; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2473 = 5'hd == _T_268[4:0] ? io_in_13_Re : _GEN_2472; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2474 = 5'he == _T_268[4:0] ? io_in_14_Re : _GEN_2473; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2475 = 5'hf == _T_268[4:0] ? io_in_15_Re : _GEN_2474; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2476 = 5'h10 == _T_268[4:0] ? io_in_16_Re : _GEN_2475; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2477 = 5'h11 == _T_268[4:0] ? io_in_17_Re : _GEN_2476; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2478 = 5'h12 == _T_268[4:0] ? io_in_18_Re : _GEN_2477; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2479 = 5'h13 == _T_268[4:0] ? io_in_19_Re : _GEN_2478; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2480 = 5'h14 == _T_268[4:0] ? io_in_20_Re : _GEN_2479; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2481 = 5'h15 == _T_268[4:0] ? io_in_21_Re : _GEN_2480; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2482 = 5'h16 == _T_268[4:0] ? io_in_22_Re : _GEN_2481; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2483 = 5'h17 == _T_268[4:0] ? io_in_23_Re : _GEN_2482; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2484 = 5'h18 == _T_268[4:0] ? io_in_24_Re : _GEN_2483; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2485 = 5'h19 == _T_268[4:0] ? io_in_25_Re : _GEN_2484; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_280 = _T_2 + 37'h17; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2497 = 5'ha == _T_280[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2498 = 5'hb == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2497; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2499 = 5'hc == _T_280[4:0] ? 32'h3f800000 : _GEN_2498; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2500 = 5'hd == _T_280[4:0] ? 32'h3f441b7c : _GEN_2499; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2501 = 5'he == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2500; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2502 = 5'hf == _T_280[4:0] ? 32'h3f800000 : _GEN_2501; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2503 = 5'h10 == _T_280[4:0] ? 32'h3f441b7c : _GEN_2502; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2504 = 5'h11 == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2503; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2505 = 5'h12 == _T_280[4:0] ? 32'h3f800000 : _GEN_2504; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2506 = 5'h13 == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2505; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2507 = 5'h14 == _T_280[4:0] ? 32'hbf708fb2 : _GEN_2506; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2508 = 5'h15 == _T_280[4:0] ? 32'h3f800000 : _GEN_2507; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2509 = 5'h16 == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2508; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2510 = 5'h17 == _T_280[4:0] ? 32'hbf708fb2 : _GEN_2509; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2511 = 5'h18 == _T_280[4:0] ? 32'h3f800000 : _GEN_2510; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2512 = 5'h19 == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2511; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2524 = 5'ha == _T_280[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2525 = 5'hb == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2524; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2526 = 5'hc == _T_280[4:0] ? 32'h80800000 : _GEN_2525; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2527 = 5'hd == _T_280[4:0] ? 32'hbf248dba : _GEN_2526; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2528 = 5'he == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2527; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2529 = 5'hf == _T_280[4:0] ? 32'h80800000 : _GEN_2528; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2530 = 5'h10 == _T_280[4:0] ? 32'hbf248dba : _GEN_2529; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2531 = 5'h11 == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2530; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2532 = 5'h12 == _T_280[4:0] ? 32'h80800000 : _GEN_2531; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2533 = 5'h13 == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2532; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2534 = 5'h14 == _T_280[4:0] ? 32'hbeaf1d40 : _GEN_2533; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2535 = 5'h15 == _T_280[4:0] ? 32'h80800000 : _GEN_2534; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2536 = 5'h16 == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2535; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2537 = 5'h17 == _T_280[4:0] ? 32'hbeaf1d40 : _GEN_2536; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2538 = 5'h18 == _T_280[4:0] ? 32'h80800000 : _GEN_2537; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2539 = 5'h19 == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2538; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2542 = 5'h1 == _T_280[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2543 = 5'h2 == _T_280[4:0] ? io_in_2_Im : _GEN_2542; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2544 = 5'h3 == _T_280[4:0] ? io_in_3_Im : _GEN_2543; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2545 = 5'h4 == _T_280[4:0] ? io_in_4_Im : _GEN_2544; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2546 = 5'h5 == _T_280[4:0] ? io_in_5_Im : _GEN_2545; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2547 = 5'h6 == _T_280[4:0] ? io_in_6_Im : _GEN_2546; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2548 = 5'h7 == _T_280[4:0] ? io_in_7_Im : _GEN_2547; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2549 = 5'h8 == _T_280[4:0] ? io_in_8_Im : _GEN_2548; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2550 = 5'h9 == _T_280[4:0] ? io_in_9_Im : _GEN_2549; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2551 = 5'ha == _T_280[4:0] ? io_in_10_Im : _GEN_2550; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2552 = 5'hb == _T_280[4:0] ? io_in_11_Im : _GEN_2551; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2553 = 5'hc == _T_280[4:0] ? io_in_12_Im : _GEN_2552; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2554 = 5'hd == _T_280[4:0] ? io_in_13_Im : _GEN_2553; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2555 = 5'he == _T_280[4:0] ? io_in_14_Im : _GEN_2554; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2556 = 5'hf == _T_280[4:0] ? io_in_15_Im : _GEN_2555; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2557 = 5'h10 == _T_280[4:0] ? io_in_16_Im : _GEN_2556; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2558 = 5'h11 == _T_280[4:0] ? io_in_17_Im : _GEN_2557; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2559 = 5'h12 == _T_280[4:0] ? io_in_18_Im : _GEN_2558; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2560 = 5'h13 == _T_280[4:0] ? io_in_19_Im : _GEN_2559; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2561 = 5'h14 == _T_280[4:0] ? io_in_20_Im : _GEN_2560; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2562 = 5'h15 == _T_280[4:0] ? io_in_21_Im : _GEN_2561; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2563 = 5'h16 == _T_280[4:0] ? io_in_22_Im : _GEN_2562; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2564 = 5'h17 == _T_280[4:0] ? io_in_23_Im : _GEN_2563; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2565 = 5'h18 == _T_280[4:0] ? io_in_24_Im : _GEN_2564; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2566 = 5'h19 == _T_280[4:0] ? io_in_25_Im : _GEN_2565; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2569 = 5'h1 == _T_280[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2570 = 5'h2 == _T_280[4:0] ? io_in_2_Re : _GEN_2569; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2571 = 5'h3 == _T_280[4:0] ? io_in_3_Re : _GEN_2570; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2572 = 5'h4 == _T_280[4:0] ? io_in_4_Re : _GEN_2571; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2573 = 5'h5 == _T_280[4:0] ? io_in_5_Re : _GEN_2572; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2574 = 5'h6 == _T_280[4:0] ? io_in_6_Re : _GEN_2573; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2575 = 5'h7 == _T_280[4:0] ? io_in_7_Re : _GEN_2574; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2576 = 5'h8 == _T_280[4:0] ? io_in_8_Re : _GEN_2575; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2577 = 5'h9 == _T_280[4:0] ? io_in_9_Re : _GEN_2576; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2578 = 5'ha == _T_280[4:0] ? io_in_10_Re : _GEN_2577; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2579 = 5'hb == _T_280[4:0] ? io_in_11_Re : _GEN_2578; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2580 = 5'hc == _T_280[4:0] ? io_in_12_Re : _GEN_2579; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2581 = 5'hd == _T_280[4:0] ? io_in_13_Re : _GEN_2580; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2582 = 5'he == _T_280[4:0] ? io_in_14_Re : _GEN_2581; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2583 = 5'hf == _T_280[4:0] ? io_in_15_Re : _GEN_2582; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2584 = 5'h10 == _T_280[4:0] ? io_in_16_Re : _GEN_2583; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2585 = 5'h11 == _T_280[4:0] ? io_in_17_Re : _GEN_2584; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2586 = 5'h12 == _T_280[4:0] ? io_in_18_Re : _GEN_2585; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2587 = 5'h13 == _T_280[4:0] ? io_in_19_Re : _GEN_2586; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2588 = 5'h14 == _T_280[4:0] ? io_in_20_Re : _GEN_2587; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2589 = 5'h15 == _T_280[4:0] ? io_in_21_Re : _GEN_2588; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2590 = 5'h16 == _T_280[4:0] ? io_in_22_Re : _GEN_2589; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2591 = 5'h17 == _T_280[4:0] ? io_in_23_Re : _GEN_2590; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2592 = 5'h18 == _T_280[4:0] ? io_in_24_Re : _GEN_2591; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2593 = 5'h19 == _T_280[4:0] ? io_in_25_Re : _GEN_2592; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_292 = _T_2 + 37'h18; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2605 = 5'ha == _T_292[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2606 = 5'hb == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2605; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2607 = 5'hc == _T_292[4:0] ? 32'h3f800000 : _GEN_2606; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2608 = 5'hd == _T_292[4:0] ? 32'h3f441b7c : _GEN_2607; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2609 = 5'he == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2608; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2610 = 5'hf == _T_292[4:0] ? 32'h3f800000 : _GEN_2609; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2611 = 5'h10 == _T_292[4:0] ? 32'h3f441b7c : _GEN_2610; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2612 = 5'h11 == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2611; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2613 = 5'h12 == _T_292[4:0] ? 32'h3f800000 : _GEN_2612; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2614 = 5'h13 == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2613; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2615 = 5'h14 == _T_292[4:0] ? 32'hbf708fb2 : _GEN_2614; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2616 = 5'h15 == _T_292[4:0] ? 32'h3f800000 : _GEN_2615; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2617 = 5'h16 == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2616; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2618 = 5'h17 == _T_292[4:0] ? 32'hbf708fb2 : _GEN_2617; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2619 = 5'h18 == _T_292[4:0] ? 32'h3f800000 : _GEN_2618; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2620 = 5'h19 == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2619; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2632 = 5'ha == _T_292[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2633 = 5'hb == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2632; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2634 = 5'hc == _T_292[4:0] ? 32'h80800000 : _GEN_2633; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2635 = 5'hd == _T_292[4:0] ? 32'hbf248dba : _GEN_2634; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2636 = 5'he == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2635; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2637 = 5'hf == _T_292[4:0] ? 32'h80800000 : _GEN_2636; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2638 = 5'h10 == _T_292[4:0] ? 32'hbf248dba : _GEN_2637; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2639 = 5'h11 == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2638; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2640 = 5'h12 == _T_292[4:0] ? 32'h80800000 : _GEN_2639; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2641 = 5'h13 == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2640; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2642 = 5'h14 == _T_292[4:0] ? 32'hbeaf1d40 : _GEN_2641; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2643 = 5'h15 == _T_292[4:0] ? 32'h80800000 : _GEN_2642; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2644 = 5'h16 == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2643; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2645 = 5'h17 == _T_292[4:0] ? 32'hbeaf1d40 : _GEN_2644; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2646 = 5'h18 == _T_292[4:0] ? 32'h80800000 : _GEN_2645; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2647 = 5'h19 == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2646; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2650 = 5'h1 == _T_292[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2651 = 5'h2 == _T_292[4:0] ? io_in_2_Im : _GEN_2650; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2652 = 5'h3 == _T_292[4:0] ? io_in_3_Im : _GEN_2651; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2653 = 5'h4 == _T_292[4:0] ? io_in_4_Im : _GEN_2652; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2654 = 5'h5 == _T_292[4:0] ? io_in_5_Im : _GEN_2653; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2655 = 5'h6 == _T_292[4:0] ? io_in_6_Im : _GEN_2654; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2656 = 5'h7 == _T_292[4:0] ? io_in_7_Im : _GEN_2655; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2657 = 5'h8 == _T_292[4:0] ? io_in_8_Im : _GEN_2656; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2658 = 5'h9 == _T_292[4:0] ? io_in_9_Im : _GEN_2657; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2659 = 5'ha == _T_292[4:0] ? io_in_10_Im : _GEN_2658; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2660 = 5'hb == _T_292[4:0] ? io_in_11_Im : _GEN_2659; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2661 = 5'hc == _T_292[4:0] ? io_in_12_Im : _GEN_2660; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2662 = 5'hd == _T_292[4:0] ? io_in_13_Im : _GEN_2661; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2663 = 5'he == _T_292[4:0] ? io_in_14_Im : _GEN_2662; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2664 = 5'hf == _T_292[4:0] ? io_in_15_Im : _GEN_2663; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2665 = 5'h10 == _T_292[4:0] ? io_in_16_Im : _GEN_2664; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2666 = 5'h11 == _T_292[4:0] ? io_in_17_Im : _GEN_2665; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2667 = 5'h12 == _T_292[4:0] ? io_in_18_Im : _GEN_2666; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2668 = 5'h13 == _T_292[4:0] ? io_in_19_Im : _GEN_2667; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2669 = 5'h14 == _T_292[4:0] ? io_in_20_Im : _GEN_2668; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2670 = 5'h15 == _T_292[4:0] ? io_in_21_Im : _GEN_2669; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2671 = 5'h16 == _T_292[4:0] ? io_in_22_Im : _GEN_2670; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2672 = 5'h17 == _T_292[4:0] ? io_in_23_Im : _GEN_2671; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2673 = 5'h18 == _T_292[4:0] ? io_in_24_Im : _GEN_2672; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2674 = 5'h19 == _T_292[4:0] ? io_in_25_Im : _GEN_2673; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2677 = 5'h1 == _T_292[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2678 = 5'h2 == _T_292[4:0] ? io_in_2_Re : _GEN_2677; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2679 = 5'h3 == _T_292[4:0] ? io_in_3_Re : _GEN_2678; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2680 = 5'h4 == _T_292[4:0] ? io_in_4_Re : _GEN_2679; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2681 = 5'h5 == _T_292[4:0] ? io_in_5_Re : _GEN_2680; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2682 = 5'h6 == _T_292[4:0] ? io_in_6_Re : _GEN_2681; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2683 = 5'h7 == _T_292[4:0] ? io_in_7_Re : _GEN_2682; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2684 = 5'h8 == _T_292[4:0] ? io_in_8_Re : _GEN_2683; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2685 = 5'h9 == _T_292[4:0] ? io_in_9_Re : _GEN_2684; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2686 = 5'ha == _T_292[4:0] ? io_in_10_Re : _GEN_2685; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2687 = 5'hb == _T_292[4:0] ? io_in_11_Re : _GEN_2686; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2688 = 5'hc == _T_292[4:0] ? io_in_12_Re : _GEN_2687; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2689 = 5'hd == _T_292[4:0] ? io_in_13_Re : _GEN_2688; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2690 = 5'he == _T_292[4:0] ? io_in_14_Re : _GEN_2689; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2691 = 5'hf == _T_292[4:0] ? io_in_15_Re : _GEN_2690; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2692 = 5'h10 == _T_292[4:0] ? io_in_16_Re : _GEN_2691; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2693 = 5'h11 == _T_292[4:0] ? io_in_17_Re : _GEN_2692; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2694 = 5'h12 == _T_292[4:0] ? io_in_18_Re : _GEN_2693; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2695 = 5'h13 == _T_292[4:0] ? io_in_19_Re : _GEN_2694; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2696 = 5'h14 == _T_292[4:0] ? io_in_20_Re : _GEN_2695; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2697 = 5'h15 == _T_292[4:0] ? io_in_21_Re : _GEN_2696; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2698 = 5'h16 == _T_292[4:0] ? io_in_22_Re : _GEN_2697; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2699 = 5'h17 == _T_292[4:0] ? io_in_23_Re : _GEN_2698; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2700 = 5'h18 == _T_292[4:0] ? io_in_24_Re : _GEN_2699; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2701 = 5'h19 == _T_292[4:0] ? io_in_25_Re : _GEN_2700; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_304 = _T_2 + 37'h19; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2713 = 5'ha == _T_304[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2714 = 5'hb == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2713; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2715 = 5'hc == _T_304[4:0] ? 32'h3f800000 : _GEN_2714; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2716 = 5'hd == _T_304[4:0] ? 32'h3f441b7c : _GEN_2715; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2717 = 5'he == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2716; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2718 = 5'hf == _T_304[4:0] ? 32'h3f800000 : _GEN_2717; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2719 = 5'h10 == _T_304[4:0] ? 32'h3f441b7c : _GEN_2718; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2720 = 5'h11 == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2719; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2721 = 5'h12 == _T_304[4:0] ? 32'h3f800000 : _GEN_2720; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2722 = 5'h13 == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2721; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2723 = 5'h14 == _T_304[4:0] ? 32'hbf708fb2 : _GEN_2722; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2724 = 5'h15 == _T_304[4:0] ? 32'h3f800000 : _GEN_2723; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2725 = 5'h16 == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2724; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2726 = 5'h17 == _T_304[4:0] ? 32'hbf708fb2 : _GEN_2725; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2727 = 5'h18 == _T_304[4:0] ? 32'h3f800000 : _GEN_2726; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2728 = 5'h19 == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2727; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2740 = 5'ha == _T_304[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2741 = 5'hb == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2740; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2742 = 5'hc == _T_304[4:0] ? 32'h80800000 : _GEN_2741; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2743 = 5'hd == _T_304[4:0] ? 32'hbf248dba : _GEN_2742; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2744 = 5'he == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2743; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2745 = 5'hf == _T_304[4:0] ? 32'h80800000 : _GEN_2744; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2746 = 5'h10 == _T_304[4:0] ? 32'hbf248dba : _GEN_2745; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2747 = 5'h11 == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2746; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2748 = 5'h12 == _T_304[4:0] ? 32'h80800000 : _GEN_2747; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2749 = 5'h13 == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2748; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2750 = 5'h14 == _T_304[4:0] ? 32'hbeaf1d40 : _GEN_2749; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2751 = 5'h15 == _T_304[4:0] ? 32'h80800000 : _GEN_2750; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2752 = 5'h16 == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2751; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2753 = 5'h17 == _T_304[4:0] ? 32'hbeaf1d40 : _GEN_2752; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2754 = 5'h18 == _T_304[4:0] ? 32'h80800000 : _GEN_2753; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2755 = 5'h19 == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2754; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2758 = 5'h1 == _T_304[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2759 = 5'h2 == _T_304[4:0] ? io_in_2_Im : _GEN_2758; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2760 = 5'h3 == _T_304[4:0] ? io_in_3_Im : _GEN_2759; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2761 = 5'h4 == _T_304[4:0] ? io_in_4_Im : _GEN_2760; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2762 = 5'h5 == _T_304[4:0] ? io_in_5_Im : _GEN_2761; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2763 = 5'h6 == _T_304[4:0] ? io_in_6_Im : _GEN_2762; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2764 = 5'h7 == _T_304[4:0] ? io_in_7_Im : _GEN_2763; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2765 = 5'h8 == _T_304[4:0] ? io_in_8_Im : _GEN_2764; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2766 = 5'h9 == _T_304[4:0] ? io_in_9_Im : _GEN_2765; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2767 = 5'ha == _T_304[4:0] ? io_in_10_Im : _GEN_2766; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2768 = 5'hb == _T_304[4:0] ? io_in_11_Im : _GEN_2767; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2769 = 5'hc == _T_304[4:0] ? io_in_12_Im : _GEN_2768; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2770 = 5'hd == _T_304[4:0] ? io_in_13_Im : _GEN_2769; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2771 = 5'he == _T_304[4:0] ? io_in_14_Im : _GEN_2770; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2772 = 5'hf == _T_304[4:0] ? io_in_15_Im : _GEN_2771; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2773 = 5'h10 == _T_304[4:0] ? io_in_16_Im : _GEN_2772; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2774 = 5'h11 == _T_304[4:0] ? io_in_17_Im : _GEN_2773; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2775 = 5'h12 == _T_304[4:0] ? io_in_18_Im : _GEN_2774; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2776 = 5'h13 == _T_304[4:0] ? io_in_19_Im : _GEN_2775; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2777 = 5'h14 == _T_304[4:0] ? io_in_20_Im : _GEN_2776; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2778 = 5'h15 == _T_304[4:0] ? io_in_21_Im : _GEN_2777; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2779 = 5'h16 == _T_304[4:0] ? io_in_22_Im : _GEN_2778; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2780 = 5'h17 == _T_304[4:0] ? io_in_23_Im : _GEN_2779; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2781 = 5'h18 == _T_304[4:0] ? io_in_24_Im : _GEN_2780; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2782 = 5'h19 == _T_304[4:0] ? io_in_25_Im : _GEN_2781; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2785 = 5'h1 == _T_304[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2786 = 5'h2 == _T_304[4:0] ? io_in_2_Re : _GEN_2785; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2787 = 5'h3 == _T_304[4:0] ? io_in_3_Re : _GEN_2786; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2788 = 5'h4 == _T_304[4:0] ? io_in_4_Re : _GEN_2787; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2789 = 5'h5 == _T_304[4:0] ? io_in_5_Re : _GEN_2788; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2790 = 5'h6 == _T_304[4:0] ? io_in_6_Re : _GEN_2789; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2791 = 5'h7 == _T_304[4:0] ? io_in_7_Re : _GEN_2790; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2792 = 5'h8 == _T_304[4:0] ? io_in_8_Re : _GEN_2791; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2793 = 5'h9 == _T_304[4:0] ? io_in_9_Re : _GEN_2792; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2794 = 5'ha == _T_304[4:0] ? io_in_10_Re : _GEN_2793; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2795 = 5'hb == _T_304[4:0] ? io_in_11_Re : _GEN_2794; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2796 = 5'hc == _T_304[4:0] ? io_in_12_Re : _GEN_2795; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2797 = 5'hd == _T_304[4:0] ? io_in_13_Re : _GEN_2796; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2798 = 5'he == _T_304[4:0] ? io_in_14_Re : _GEN_2797; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2799 = 5'hf == _T_304[4:0] ? io_in_15_Re : _GEN_2798; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2800 = 5'h10 == _T_304[4:0] ? io_in_16_Re : _GEN_2799; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2801 = 5'h11 == _T_304[4:0] ? io_in_17_Re : _GEN_2800; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2802 = 5'h12 == _T_304[4:0] ? io_in_18_Re : _GEN_2801; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2803 = 5'h13 == _T_304[4:0] ? io_in_19_Re : _GEN_2802; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2804 = 5'h14 == _T_304[4:0] ? io_in_20_Re : _GEN_2803; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2805 = 5'h15 == _T_304[4:0] ? io_in_21_Re : _GEN_2804; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2806 = 5'h16 == _T_304[4:0] ? io_in_22_Re : _GEN_2805; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2807 = 5'h17 == _T_304[4:0] ? io_in_23_Re : _GEN_2806; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2808 = 5'h18 == _T_304[4:0] ? io_in_24_Re : _GEN_2807; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2809 = 5'h19 == _T_304[4:0] ? io_in_25_Re : _GEN_2808; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_316 = _T_2 + 37'h1a; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2821 = 5'ha == _T_316[4:0] ? 32'h3f441b7c : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2822 = 5'hb == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2821; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2823 = 5'hc == _T_316[4:0] ? 32'h3f800000 : _GEN_2822; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2824 = 5'hd == _T_316[4:0] ? 32'h3f441b7c : _GEN_2823; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2825 = 5'he == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2824; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2826 = 5'hf == _T_316[4:0] ? 32'h3f800000 : _GEN_2825; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2827 = 5'h10 == _T_316[4:0] ? 32'h3f441b7c : _GEN_2826; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2828 = 5'h11 == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2827; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2829 = 5'h12 == _T_316[4:0] ? 32'h3f800000 : _GEN_2828; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2830 = 5'h13 == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2829; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2831 = 5'h14 == _T_316[4:0] ? 32'hbf708fb2 : _GEN_2830; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2832 = 5'h15 == _T_316[4:0] ? 32'h3f800000 : _GEN_2831; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2833 = 5'h16 == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2832; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2834 = 5'h17 == _T_316[4:0] ? 32'hbf708fb2 : _GEN_2833; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2835 = 5'h18 == _T_316[4:0] ? 32'h3f800000 : _GEN_2834; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2836 = 5'h19 == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2835; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2848 = 5'ha == _T_316[4:0] ? 32'hbf248dba : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2849 = 5'hb == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2848; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2850 = 5'hc == _T_316[4:0] ? 32'h80800000 : _GEN_2849; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2851 = 5'hd == _T_316[4:0] ? 32'hbf248dba : _GEN_2850; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2852 = 5'he == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2851; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2853 = 5'hf == _T_316[4:0] ? 32'h80800000 : _GEN_2852; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2854 = 5'h10 == _T_316[4:0] ? 32'hbf248dba : _GEN_2853; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2855 = 5'h11 == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2854; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2856 = 5'h12 == _T_316[4:0] ? 32'h80800000 : _GEN_2855; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2857 = 5'h13 == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2856; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2858 = 5'h14 == _T_316[4:0] ? 32'hbeaf1d40 : _GEN_2857; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2859 = 5'h15 == _T_316[4:0] ? 32'h80800000 : _GEN_2858; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2860 = 5'h16 == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2859; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2861 = 5'h17 == _T_316[4:0] ? 32'hbeaf1d40 : _GEN_2860; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2862 = 5'h18 == _T_316[4:0] ? 32'h80800000 : _GEN_2861; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2863 = 5'h19 == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2862; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2866 = 5'h1 == _T_316[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2867 = 5'h2 == _T_316[4:0] ? io_in_2_Im : _GEN_2866; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2868 = 5'h3 == _T_316[4:0] ? io_in_3_Im : _GEN_2867; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2869 = 5'h4 == _T_316[4:0] ? io_in_4_Im : _GEN_2868; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2870 = 5'h5 == _T_316[4:0] ? io_in_5_Im : _GEN_2869; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2871 = 5'h6 == _T_316[4:0] ? io_in_6_Im : _GEN_2870; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2872 = 5'h7 == _T_316[4:0] ? io_in_7_Im : _GEN_2871; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2873 = 5'h8 == _T_316[4:0] ? io_in_8_Im : _GEN_2872; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2874 = 5'h9 == _T_316[4:0] ? io_in_9_Im : _GEN_2873; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2875 = 5'ha == _T_316[4:0] ? io_in_10_Im : _GEN_2874; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2876 = 5'hb == _T_316[4:0] ? io_in_11_Im : _GEN_2875; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2877 = 5'hc == _T_316[4:0] ? io_in_12_Im : _GEN_2876; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2878 = 5'hd == _T_316[4:0] ? io_in_13_Im : _GEN_2877; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2879 = 5'he == _T_316[4:0] ? io_in_14_Im : _GEN_2878; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2880 = 5'hf == _T_316[4:0] ? io_in_15_Im : _GEN_2879; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2881 = 5'h10 == _T_316[4:0] ? io_in_16_Im : _GEN_2880; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2882 = 5'h11 == _T_316[4:0] ? io_in_17_Im : _GEN_2881; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2883 = 5'h12 == _T_316[4:0] ? io_in_18_Im : _GEN_2882; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2884 = 5'h13 == _T_316[4:0] ? io_in_19_Im : _GEN_2883; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2885 = 5'h14 == _T_316[4:0] ? io_in_20_Im : _GEN_2884; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2886 = 5'h15 == _T_316[4:0] ? io_in_21_Im : _GEN_2885; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2887 = 5'h16 == _T_316[4:0] ? io_in_22_Im : _GEN_2886; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2888 = 5'h17 == _T_316[4:0] ? io_in_23_Im : _GEN_2887; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2889 = 5'h18 == _T_316[4:0] ? io_in_24_Im : _GEN_2888; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2890 = 5'h19 == _T_316[4:0] ? io_in_25_Im : _GEN_2889; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2893 = 5'h1 == _T_316[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2894 = 5'h2 == _T_316[4:0] ? io_in_2_Re : _GEN_2893; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2895 = 5'h3 == _T_316[4:0] ? io_in_3_Re : _GEN_2894; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2896 = 5'h4 == _T_316[4:0] ? io_in_4_Re : _GEN_2895; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2897 = 5'h5 == _T_316[4:0] ? io_in_5_Re : _GEN_2896; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2898 = 5'h6 == _T_316[4:0] ? io_in_6_Re : _GEN_2897; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2899 = 5'h7 == _T_316[4:0] ? io_in_7_Re : _GEN_2898; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2900 = 5'h8 == _T_316[4:0] ? io_in_8_Re : _GEN_2899; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2901 = 5'h9 == _T_316[4:0] ? io_in_9_Re : _GEN_2900; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2902 = 5'ha == _T_316[4:0] ? io_in_10_Re : _GEN_2901; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2903 = 5'hb == _T_316[4:0] ? io_in_11_Re : _GEN_2902; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2904 = 5'hc == _T_316[4:0] ? io_in_12_Re : _GEN_2903; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2905 = 5'hd == _T_316[4:0] ? io_in_13_Re : _GEN_2904; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2906 = 5'he == _T_316[4:0] ? io_in_14_Re : _GEN_2905; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2907 = 5'hf == _T_316[4:0] ? io_in_15_Re : _GEN_2906; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2908 = 5'h10 == _T_316[4:0] ? io_in_16_Re : _GEN_2907; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2909 = 5'h11 == _T_316[4:0] ? io_in_17_Re : _GEN_2908; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2910 = 5'h12 == _T_316[4:0] ? io_in_18_Re : _GEN_2909; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2911 = 5'h13 == _T_316[4:0] ? io_in_19_Re : _GEN_2910; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2912 = 5'h14 == _T_316[4:0] ? io_in_20_Re : _GEN_2911; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2913 = 5'h15 == _T_316[4:0] ? io_in_21_Re : _GEN_2912; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2914 = 5'h16 == _T_316[4:0] ? io_in_22_Re : _GEN_2913; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2915 = 5'h17 == _T_316[4:0] ? io_in_23_Re : _GEN_2914; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2916 = 5'h18 == _T_316[4:0] ? io_in_24_Re : _GEN_2915; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2917 = 5'h19 == _T_316[4:0] ? io_in_25_Re : _GEN_2916; // @[FFTDesigns.scala 543:{23,23}]
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_clock),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_1_clock),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_2_clock),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_3_clock),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_4_clock),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_5_clock),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_6_clock),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_7_clock),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_8_clock),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_9_clock),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_10_clock),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_11_clock),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_12 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_12_clock),
    .io_in_a_Re(FPComplexMult_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_12_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_13 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_13_clock),
    .io_in_a_Re(FPComplexMult_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_13_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_14 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_14_clock),
    .io_in_a_Re(FPComplexMult_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_14_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_15 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_15_clock),
    .io_in_a_Re(FPComplexMult_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_15_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_16 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_16_clock),
    .io_in_a_Re(FPComplexMult_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_16_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_16_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_16_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_16_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_17 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_17_clock),
    .io_in_a_Re(FPComplexMult_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_17_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_17_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_17_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_17_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_18 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_18_clock),
    .io_in_a_Re(FPComplexMult_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_18_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_18_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_18_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_18_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_19 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_19_clock),
    .io_in_a_Re(FPComplexMult_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_19_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_19_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_19_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_19_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_20 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_20_clock),
    .io_in_a_Re(FPComplexMult_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_20_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_20_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_20_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_20_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_21 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_21_clock),
    .io_in_a_Re(FPComplexMult_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_21_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_21_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_21_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_21_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_22 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_22_clock),
    .io_in_a_Re(FPComplexMult_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_22_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_22_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_22_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_22_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_23 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_23_clock),
    .io_in_a_Re(FPComplexMult_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_23_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_23_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_23_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_23_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_24 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_24_clock),
    .io_in_a_Re(FPComplexMult_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_24_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_24_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_24_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_24_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_25 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_25_clock),
    .io_in_a_Re(FPComplexMult_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_25_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_25_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_25_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_25_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_26 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_26_clock),
    .io_in_a_Re(FPComplexMult_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_26_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_26_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_26_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_26_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_12_Re = FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_12_Im = FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_13_Re = FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_13_Im = FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_14_Re = FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_14_Im = FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_15_Re = FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_15_Im = FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_16_Re = FPComplexMult_16_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_16_Im = FPComplexMult_16_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_17_Re = FPComplexMult_17_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_17_Im = FPComplexMult_17_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_18_Re = FPComplexMult_18_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_18_Im = FPComplexMult_18_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_19_Re = FPComplexMult_19_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_19_Im = FPComplexMult_19_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_20_Re = FPComplexMult_20_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_20_Im = FPComplexMult_20_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_21_Re = FPComplexMult_21_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_21_Im = FPComplexMult_21_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_22_Re = FPComplexMult_22_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_22_Im = FPComplexMult_22_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_23_Re = FPComplexMult_23_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_23_Im = FPComplexMult_23_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_24_Re = FPComplexMult_24_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_24_Im = FPComplexMult_24_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_25_Re = FPComplexMult_25_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_25_Im = FPComplexMult_25_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_26_Re = FPComplexMult_26_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_26_Im = FPComplexMult_26_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_io_in_a_Re = 5'h1a == _T_3[4:0] ? 32'hbf708fb2 : _GEN_28; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_io_in_a_Im = 5'h1a == _T_3[4:0] ? 32'hbeaf1d40 : _GEN_55; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_io_in_b_Re = 5'h1a == _T_3[4:0] ? io_in_26_Re : _GEN_109; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_io_in_b_Im = 5'h1a == _T_3[4:0] ? io_in_26_Im : _GEN_82; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_io_in_a_Re = 5'h1a == _T_16[4:0] ? 32'hbf708fb2 : _GEN_136; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_1_io_in_a_Im = 5'h1a == _T_16[4:0] ? 32'hbeaf1d40 : _GEN_163; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_1_io_in_b_Re = 5'h1a == _T_16[4:0] ? io_in_26_Re : _GEN_217; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_1_io_in_b_Im = 5'h1a == _T_16[4:0] ? io_in_26_Im : _GEN_190; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_io_in_a_Re = 5'h1a == _T_28[4:0] ? 32'hbf708fb2 : _GEN_244; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_2_io_in_a_Im = 5'h1a == _T_28[4:0] ? 32'hbeaf1d40 : _GEN_271; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_2_io_in_b_Re = 5'h1a == _T_28[4:0] ? io_in_26_Re : _GEN_325; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_2_io_in_b_Im = 5'h1a == _T_28[4:0] ? io_in_26_Im : _GEN_298; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_io_in_a_Re = 5'h1a == _T_40[4:0] ? 32'hbf708fb2 : _GEN_352; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_3_io_in_a_Im = 5'h1a == _T_40[4:0] ? 32'hbeaf1d40 : _GEN_379; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_3_io_in_b_Re = 5'h1a == _T_40[4:0] ? io_in_26_Re : _GEN_433; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_3_io_in_b_Im = 5'h1a == _T_40[4:0] ? io_in_26_Im : _GEN_406; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_io_in_a_Re = 5'h1a == _T_52[4:0] ? 32'hbf708fb2 : _GEN_460; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_4_io_in_a_Im = 5'h1a == _T_52[4:0] ? 32'hbeaf1d40 : _GEN_487; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_4_io_in_b_Re = 5'h1a == _T_52[4:0] ? io_in_26_Re : _GEN_541; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_4_io_in_b_Im = 5'h1a == _T_52[4:0] ? io_in_26_Im : _GEN_514; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_io_in_a_Re = 5'h1a == _T_64[4:0] ? 32'hbf708fb2 : _GEN_568; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_5_io_in_a_Im = 5'h1a == _T_64[4:0] ? 32'hbeaf1d40 : _GEN_595; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_5_io_in_b_Re = 5'h1a == _T_64[4:0] ? io_in_26_Re : _GEN_649; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_5_io_in_b_Im = 5'h1a == _T_64[4:0] ? io_in_26_Im : _GEN_622; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_io_in_a_Re = 5'h1a == _T_76[4:0] ? 32'hbf708fb2 : _GEN_676; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_6_io_in_a_Im = 5'h1a == _T_76[4:0] ? 32'hbeaf1d40 : _GEN_703; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_6_io_in_b_Re = 5'h1a == _T_76[4:0] ? io_in_26_Re : _GEN_757; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_6_io_in_b_Im = 5'h1a == _T_76[4:0] ? io_in_26_Im : _GEN_730; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_io_in_a_Re = 5'h1a == _T_88[4:0] ? 32'hbf708fb2 : _GEN_784; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_7_io_in_a_Im = 5'h1a == _T_88[4:0] ? 32'hbeaf1d40 : _GEN_811; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_7_io_in_b_Re = 5'h1a == _T_88[4:0] ? io_in_26_Re : _GEN_865; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_7_io_in_b_Im = 5'h1a == _T_88[4:0] ? io_in_26_Im : _GEN_838; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_io_in_a_Re = 5'h1a == _T_100[4:0] ? 32'hbf708fb2 : _GEN_892; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_8_io_in_a_Im = 5'h1a == _T_100[4:0] ? 32'hbeaf1d40 : _GEN_919; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_8_io_in_b_Re = 5'h1a == _T_100[4:0] ? io_in_26_Re : _GEN_973; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_8_io_in_b_Im = 5'h1a == _T_100[4:0] ? io_in_26_Im : _GEN_946; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_io_in_a_Re = 5'h1a == _T_112[4:0] ? 32'hbf708fb2 : _GEN_1000; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_9_io_in_a_Im = 5'h1a == _T_112[4:0] ? 32'hbeaf1d40 : _GEN_1027; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_9_io_in_b_Re = 5'h1a == _T_112[4:0] ? io_in_26_Re : _GEN_1081; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_9_io_in_b_Im = 5'h1a == _T_112[4:0] ? io_in_26_Im : _GEN_1054; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_io_in_a_Re = 5'h1a == _T_124[4:0] ? 32'hbf708fb2 : _GEN_1108; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_10_io_in_a_Im = 5'h1a == _T_124[4:0] ? 32'hbeaf1d40 : _GEN_1135; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_10_io_in_b_Re = 5'h1a == _T_124[4:0] ? io_in_26_Re : _GEN_1189; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_10_io_in_b_Im = 5'h1a == _T_124[4:0] ? io_in_26_Im : _GEN_1162; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_io_in_a_Re = 5'h1a == _T_136[4:0] ? 32'hbf708fb2 : _GEN_1216; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_11_io_in_a_Im = 5'h1a == _T_136[4:0] ? 32'hbeaf1d40 : _GEN_1243; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_11_io_in_b_Re = 5'h1a == _T_136[4:0] ? io_in_26_Re : _GEN_1297; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_11_io_in_b_Im = 5'h1a == _T_136[4:0] ? io_in_26_Im : _GEN_1270; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_12_clock = clock;
  assign FPComplexMult_12_io_in_a_Re = 5'h1a == _T_148[4:0] ? 32'hbf708fb2 : _GEN_1324; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_12_io_in_a_Im = 5'h1a == _T_148[4:0] ? 32'hbeaf1d40 : _GEN_1351; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_12_io_in_b_Re = 5'h1a == _T_148[4:0] ? io_in_26_Re : _GEN_1405; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_12_io_in_b_Im = 5'h1a == _T_148[4:0] ? io_in_26_Im : _GEN_1378; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_13_clock = clock;
  assign FPComplexMult_13_io_in_a_Re = 5'h1a == _T_160[4:0] ? 32'hbf708fb2 : _GEN_1432; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_13_io_in_a_Im = 5'h1a == _T_160[4:0] ? 32'hbeaf1d40 : _GEN_1459; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_13_io_in_b_Re = 5'h1a == _T_160[4:0] ? io_in_26_Re : _GEN_1513; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_13_io_in_b_Im = 5'h1a == _T_160[4:0] ? io_in_26_Im : _GEN_1486; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_14_clock = clock;
  assign FPComplexMult_14_io_in_a_Re = 5'h1a == _T_172[4:0] ? 32'hbf708fb2 : _GEN_1540; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_14_io_in_a_Im = 5'h1a == _T_172[4:0] ? 32'hbeaf1d40 : _GEN_1567; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_14_io_in_b_Re = 5'h1a == _T_172[4:0] ? io_in_26_Re : _GEN_1621; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_14_io_in_b_Im = 5'h1a == _T_172[4:0] ? io_in_26_Im : _GEN_1594; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_15_clock = clock;
  assign FPComplexMult_15_io_in_a_Re = 5'h1a == _T_184[4:0] ? 32'hbf708fb2 : _GEN_1648; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_15_io_in_a_Im = 5'h1a == _T_184[4:0] ? 32'hbeaf1d40 : _GEN_1675; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_15_io_in_b_Re = 5'h1a == _T_184[4:0] ? io_in_26_Re : _GEN_1729; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_15_io_in_b_Im = 5'h1a == _T_184[4:0] ? io_in_26_Im : _GEN_1702; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_16_clock = clock;
  assign FPComplexMult_16_io_in_a_Re = 5'h1a == _T_196[4:0] ? 32'hbf708fb2 : _GEN_1756; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_16_io_in_a_Im = 5'h1a == _T_196[4:0] ? 32'hbeaf1d40 : _GEN_1783; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_16_io_in_b_Re = 5'h1a == _T_196[4:0] ? io_in_26_Re : _GEN_1837; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_16_io_in_b_Im = 5'h1a == _T_196[4:0] ? io_in_26_Im : _GEN_1810; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_17_clock = clock;
  assign FPComplexMult_17_io_in_a_Re = 5'h1a == _T_208[4:0] ? 32'hbf708fb2 : _GEN_1864; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_17_io_in_a_Im = 5'h1a == _T_208[4:0] ? 32'hbeaf1d40 : _GEN_1891; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_17_io_in_b_Re = 5'h1a == _T_208[4:0] ? io_in_26_Re : _GEN_1945; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_17_io_in_b_Im = 5'h1a == _T_208[4:0] ? io_in_26_Im : _GEN_1918; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_18_clock = clock;
  assign FPComplexMult_18_io_in_a_Re = 5'h1a == _T_220[4:0] ? 32'hbf708fb2 : _GEN_1972; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_18_io_in_a_Im = 5'h1a == _T_220[4:0] ? 32'hbeaf1d40 : _GEN_1999; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_18_io_in_b_Re = 5'h1a == _T_220[4:0] ? io_in_26_Re : _GEN_2053; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_18_io_in_b_Im = 5'h1a == _T_220[4:0] ? io_in_26_Im : _GEN_2026; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_19_clock = clock;
  assign FPComplexMult_19_io_in_a_Re = 5'h1a == _T_232[4:0] ? 32'hbf708fb2 : _GEN_2080; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_19_io_in_a_Im = 5'h1a == _T_232[4:0] ? 32'hbeaf1d40 : _GEN_2107; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_19_io_in_b_Re = 5'h1a == _T_232[4:0] ? io_in_26_Re : _GEN_2161; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_19_io_in_b_Im = 5'h1a == _T_232[4:0] ? io_in_26_Im : _GEN_2134; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_20_clock = clock;
  assign FPComplexMult_20_io_in_a_Re = 5'h1a == _T_244[4:0] ? 32'hbf708fb2 : _GEN_2188; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_20_io_in_a_Im = 5'h1a == _T_244[4:0] ? 32'hbeaf1d40 : _GEN_2215; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_20_io_in_b_Re = 5'h1a == _T_244[4:0] ? io_in_26_Re : _GEN_2269; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_20_io_in_b_Im = 5'h1a == _T_244[4:0] ? io_in_26_Im : _GEN_2242; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_21_clock = clock;
  assign FPComplexMult_21_io_in_a_Re = 5'h1a == _T_256[4:0] ? 32'hbf708fb2 : _GEN_2296; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_21_io_in_a_Im = 5'h1a == _T_256[4:0] ? 32'hbeaf1d40 : _GEN_2323; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_21_io_in_b_Re = 5'h1a == _T_256[4:0] ? io_in_26_Re : _GEN_2377; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_21_io_in_b_Im = 5'h1a == _T_256[4:0] ? io_in_26_Im : _GEN_2350; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_22_clock = clock;
  assign FPComplexMult_22_io_in_a_Re = 5'h1a == _T_268[4:0] ? 32'hbf708fb2 : _GEN_2404; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_22_io_in_a_Im = 5'h1a == _T_268[4:0] ? 32'hbeaf1d40 : _GEN_2431; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_22_io_in_b_Re = 5'h1a == _T_268[4:0] ? io_in_26_Re : _GEN_2485; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_22_io_in_b_Im = 5'h1a == _T_268[4:0] ? io_in_26_Im : _GEN_2458; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_23_clock = clock;
  assign FPComplexMult_23_io_in_a_Re = 5'h1a == _T_280[4:0] ? 32'hbf708fb2 : _GEN_2512; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_23_io_in_a_Im = 5'h1a == _T_280[4:0] ? 32'hbeaf1d40 : _GEN_2539; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_23_io_in_b_Re = 5'h1a == _T_280[4:0] ? io_in_26_Re : _GEN_2593; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_23_io_in_b_Im = 5'h1a == _T_280[4:0] ? io_in_26_Im : _GEN_2566; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_24_clock = clock;
  assign FPComplexMult_24_io_in_a_Re = 5'h1a == _T_292[4:0] ? 32'hbf708fb2 : _GEN_2620; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_24_io_in_a_Im = 5'h1a == _T_292[4:0] ? 32'hbeaf1d40 : _GEN_2647; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_24_io_in_b_Re = 5'h1a == _T_292[4:0] ? io_in_26_Re : _GEN_2701; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_24_io_in_b_Im = 5'h1a == _T_292[4:0] ? io_in_26_Im : _GEN_2674; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_25_clock = clock;
  assign FPComplexMult_25_io_in_a_Re = 5'h1a == _T_304[4:0] ? 32'hbf708fb2 : _GEN_2728; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_25_io_in_a_Im = 5'h1a == _T_304[4:0] ? 32'hbeaf1d40 : _GEN_2755; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_25_io_in_b_Re = 5'h1a == _T_304[4:0] ? io_in_26_Re : _GEN_2809; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_25_io_in_b_Im = 5'h1a == _T_304[4:0] ? io_in_26_Im : _GEN_2782; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_26_clock = clock;
  assign FPComplexMult_26_io_in_a_Re = 5'h1a == _T_316[4:0] ? 32'hbf708fb2 : _GEN_2836; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_26_io_in_a_Im = 5'h1a == _T_316[4:0] ? 32'hbeaf1d40 : _GEN_2863; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_26_io_in_b_Re = 5'h1a == _T_316[4:0] ? io_in_26_Re : _GEN_2917; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_26_io_in_b_Im = 5'h1a == _T_316[4:0] ? io_in_26_Im : _GEN_2890; // @[FFTDesigns.scala 543:{23,23}]
  always @(posedge clock) begin
    if (cnt2 == 32'h1) begin // @[FFTDesigns.scala 529:38]
      if (cnt == 32'h0) begin // @[FFTDesigns.scala 531:32]
        cnt <= 32'h0; // @[FFTDesigns.scala 532:13]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 534:13]
      end
    end
    if (cnt2 == 32'h1) begin // @[FFTDesigns.scala 529:38]
      cnt2 <= 32'h0; // @[FFTDesigns.scala 530:12]
    end else begin
      cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 538:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cnt2 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactors_1(
  input         clock,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_12_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_13_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_14_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_15_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_16_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_16_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_17_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_17_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_18_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_18_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_19_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_19_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_20_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_20_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_21_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_21_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_22_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_22_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_23_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_23_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_24_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_24_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_25_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_25_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  wire  FPComplexMult_26_clock; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_a_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_a_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_b_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_in_b_Im; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_out_s_Re; // @[FFTDesigns.scala 524:26]
  wire [31:0] FPComplexMult_26_io_out_s_Im; // @[FFTDesigns.scala 524:26]
  reg [31:0] cnt; // @[FFTDesigns.scala 527:18]
  reg [31:0] cnt2; // @[FFTDesigns.scala 528:19]
  wire [31:0] _cnt_T_1 = cnt + 32'h1; // @[FFTDesigns.scala 534:20]
  wire [31:0] _cnt2_T_1 = cnt2 + 32'h1; // @[FFTDesigns.scala 538:20]
  wire [36:0] _T_2 = cnt * 5'h1b; // @[FFTDesigns.scala 541:58]
  wire [37:0] _T_3 = {{1'd0}, _T_2}; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_7 = 5'h4 == _T_3[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_8 = 5'h5 == _T_3[4:0] ? 32'h3f64c51a : _GEN_7; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_9 = 5'h6 == _T_3[4:0] ? 32'h3f800000 : _GEN_8; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_10 = 5'h7 == _T_3[4:0] ? 32'h3f64c51a : _GEN_9; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_11 = 5'h8 == _T_3[4:0] ? 32'h3f18df62 : _GEN_10; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_12 = 5'h9 == _T_3[4:0] ? 32'h3f800000 : _GEN_11; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_13 = 5'ha == _T_3[4:0] ? 32'h3f441b7c : _GEN_12; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_14 = 5'hb == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_13; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_15 = 5'hc == _T_3[4:0] ? 32'h3f800000 : _GEN_14; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_16 = 5'hd == _T_3[4:0] ? 32'h3f18df62 : _GEN_15; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_17 = 5'he == _T_3[4:0] ? 32'hbe92d7dc : _GEN_16; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_18 = 5'hf == _T_3[4:0] ? 32'h3f800000 : _GEN_17; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_19 = 5'h10 == _T_3[4:0] ? 32'h3ecacaf4 : _GEN_18; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_20 = 5'h11 == _T_3[4:0] ? 32'hbf2fad88 : _GEN_19; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_21 = 5'h12 == _T_3[4:0] ? 32'h3f800000 : _GEN_20; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_22 = 5'h13 == _T_3[4:0] ? 32'h3e31d0d0 : _GEN_21; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_23 = 5'h14 == _T_3[4:0] ? 32'hbf708fb2 : _GEN_22; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_24 = 5'h15 == _T_3[4:0] ? 32'h3f800000 : _GEN_23; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_25 = 5'h16 == _T_3[4:0] ? 32'hbd6e2940 : _GEN_24; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_26 = 5'h17 == _T_3[4:0] ? 32'hbf7e44de : _GEN_25; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_27 = 5'h18 == _T_3[4:0] ? 32'h3f800000 : _GEN_26; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_28 = 5'h19 == _T_3[4:0] ? 32'hbe92d7dc : _GEN_27; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_34 = 5'h4 == _T_3[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_35 = 5'h5 == _T_3[4:0] ? 32'hbee5c900 : _GEN_34; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_36 = 5'h6 == _T_3[4:0] ? 32'h80800000 : _GEN_35; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_37 = 5'h7 == _T_3[4:0] ? 32'hbee5c900 : _GEN_36; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_38 = 5'h8 == _T_3[4:0] ? 32'hbf4d57f2 : _GEN_37; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_39 = 5'h9 == _T_3[4:0] ? 32'h80800000 : _GEN_38; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_40 = 5'ha == _T_3[4:0] ? 32'hbf248dba : _GEN_39; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_41 = 5'hb == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_40; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_42 = 5'hc == _T_3[4:0] ? 32'h80800000 : _GEN_41; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_43 = 5'hd == _T_3[4:0] ? 32'hbf4d57f2 : _GEN_42; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_44 = 5'he == _T_3[4:0] ? 32'hbf753ecc : _GEN_43; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_45 = 5'hf == _T_3[4:0] ? 32'h80800000 : _GEN_44; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_46 = 5'h10 == _T_3[4:0] ? 32'hbf6b1034 : _GEN_45; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_47 = 5'h11 == _T_3[4:0] ? 32'hbf3a3528 : _GEN_46; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_48 = 5'h12 == _T_3[4:0] ? 32'h80800000 : _GEN_47; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_49 = 5'h13 == _T_3[4:0] ? 32'hbf7c1c5c : _GEN_48; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_50 = 5'h14 == _T_3[4:0] ? 32'hbeaf1d40 : _GEN_49; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_51 = 5'h15 == _T_3[4:0] ? 32'h80800000 : _GEN_50; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_52 = 5'h16 == _T_3[4:0] ? 32'hbf7f911e : _GEN_51; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_53 = 5'h17 == _T_3[4:0] ? 32'h3dedc210 : _GEN_52; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_54 = 5'h18 == _T_3[4:0] ? 32'h80800000 : _GEN_53; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_55 = 5'h19 == _T_3[4:0] ? 32'hbf753ecc : _GEN_54; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_58 = 5'h1 == _T_3[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_59 = 5'h2 == _T_3[4:0] ? io_in_2_Im : _GEN_58; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_60 = 5'h3 == _T_3[4:0] ? io_in_3_Im : _GEN_59; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_61 = 5'h4 == _T_3[4:0] ? io_in_4_Im : _GEN_60; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_62 = 5'h5 == _T_3[4:0] ? io_in_5_Im : _GEN_61; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_63 = 5'h6 == _T_3[4:0] ? io_in_6_Im : _GEN_62; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_64 = 5'h7 == _T_3[4:0] ? io_in_7_Im : _GEN_63; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_65 = 5'h8 == _T_3[4:0] ? io_in_8_Im : _GEN_64; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_66 = 5'h9 == _T_3[4:0] ? io_in_9_Im : _GEN_65; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_67 = 5'ha == _T_3[4:0] ? io_in_10_Im : _GEN_66; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_68 = 5'hb == _T_3[4:0] ? io_in_11_Im : _GEN_67; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_69 = 5'hc == _T_3[4:0] ? io_in_12_Im : _GEN_68; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_70 = 5'hd == _T_3[4:0] ? io_in_13_Im : _GEN_69; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_71 = 5'he == _T_3[4:0] ? io_in_14_Im : _GEN_70; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_72 = 5'hf == _T_3[4:0] ? io_in_15_Im : _GEN_71; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_73 = 5'h10 == _T_3[4:0] ? io_in_16_Im : _GEN_72; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_74 = 5'h11 == _T_3[4:0] ? io_in_17_Im : _GEN_73; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_75 = 5'h12 == _T_3[4:0] ? io_in_18_Im : _GEN_74; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_76 = 5'h13 == _T_3[4:0] ? io_in_19_Im : _GEN_75; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_77 = 5'h14 == _T_3[4:0] ? io_in_20_Im : _GEN_76; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_78 = 5'h15 == _T_3[4:0] ? io_in_21_Im : _GEN_77; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_79 = 5'h16 == _T_3[4:0] ? io_in_22_Im : _GEN_78; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_80 = 5'h17 == _T_3[4:0] ? io_in_23_Im : _GEN_79; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_81 = 5'h18 == _T_3[4:0] ? io_in_24_Im : _GEN_80; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_82 = 5'h19 == _T_3[4:0] ? io_in_25_Im : _GEN_81; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_85 = 5'h1 == _T_3[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_86 = 5'h2 == _T_3[4:0] ? io_in_2_Re : _GEN_85; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_87 = 5'h3 == _T_3[4:0] ? io_in_3_Re : _GEN_86; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_88 = 5'h4 == _T_3[4:0] ? io_in_4_Re : _GEN_87; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_89 = 5'h5 == _T_3[4:0] ? io_in_5_Re : _GEN_88; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_90 = 5'h6 == _T_3[4:0] ? io_in_6_Re : _GEN_89; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_91 = 5'h7 == _T_3[4:0] ? io_in_7_Re : _GEN_90; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_92 = 5'h8 == _T_3[4:0] ? io_in_8_Re : _GEN_91; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_93 = 5'h9 == _T_3[4:0] ? io_in_9_Re : _GEN_92; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_94 = 5'ha == _T_3[4:0] ? io_in_10_Re : _GEN_93; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_95 = 5'hb == _T_3[4:0] ? io_in_11_Re : _GEN_94; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_96 = 5'hc == _T_3[4:0] ? io_in_12_Re : _GEN_95; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_97 = 5'hd == _T_3[4:0] ? io_in_13_Re : _GEN_96; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_98 = 5'he == _T_3[4:0] ? io_in_14_Re : _GEN_97; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_99 = 5'hf == _T_3[4:0] ? io_in_15_Re : _GEN_98; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_100 = 5'h10 == _T_3[4:0] ? io_in_16_Re : _GEN_99; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_101 = 5'h11 == _T_3[4:0] ? io_in_17_Re : _GEN_100; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_102 = 5'h12 == _T_3[4:0] ? io_in_18_Re : _GEN_101; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_103 = 5'h13 == _T_3[4:0] ? io_in_19_Re : _GEN_102; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_104 = 5'h14 == _T_3[4:0] ? io_in_20_Re : _GEN_103; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_105 = 5'h15 == _T_3[4:0] ? io_in_21_Re : _GEN_104; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_106 = 5'h16 == _T_3[4:0] ? io_in_22_Re : _GEN_105; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_107 = 5'h17 == _T_3[4:0] ? io_in_23_Re : _GEN_106; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_108 = 5'h18 == _T_3[4:0] ? io_in_24_Re : _GEN_107; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_109 = 5'h19 == _T_3[4:0] ? io_in_25_Re : _GEN_108; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_16 = _T_2 + 37'h1; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_115 = 5'h4 == _T_16[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_116 = 5'h5 == _T_16[4:0] ? 32'h3f64c51a : _GEN_115; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_117 = 5'h6 == _T_16[4:0] ? 32'h3f800000 : _GEN_116; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_118 = 5'h7 == _T_16[4:0] ? 32'h3f64c51a : _GEN_117; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_119 = 5'h8 == _T_16[4:0] ? 32'h3f18df62 : _GEN_118; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_120 = 5'h9 == _T_16[4:0] ? 32'h3f800000 : _GEN_119; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_121 = 5'ha == _T_16[4:0] ? 32'h3f441b7c : _GEN_120; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_122 = 5'hb == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_121; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_123 = 5'hc == _T_16[4:0] ? 32'h3f800000 : _GEN_122; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_124 = 5'hd == _T_16[4:0] ? 32'h3f18df62 : _GEN_123; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_125 = 5'he == _T_16[4:0] ? 32'hbe92d7dc : _GEN_124; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_126 = 5'hf == _T_16[4:0] ? 32'h3f800000 : _GEN_125; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_127 = 5'h10 == _T_16[4:0] ? 32'h3ecacaf4 : _GEN_126; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_128 = 5'h11 == _T_16[4:0] ? 32'hbf2fad88 : _GEN_127; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_129 = 5'h12 == _T_16[4:0] ? 32'h3f800000 : _GEN_128; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_130 = 5'h13 == _T_16[4:0] ? 32'h3e31d0d0 : _GEN_129; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_131 = 5'h14 == _T_16[4:0] ? 32'hbf708fb2 : _GEN_130; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_132 = 5'h15 == _T_16[4:0] ? 32'h3f800000 : _GEN_131; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_133 = 5'h16 == _T_16[4:0] ? 32'hbd6e2940 : _GEN_132; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_134 = 5'h17 == _T_16[4:0] ? 32'hbf7e44de : _GEN_133; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_135 = 5'h18 == _T_16[4:0] ? 32'h3f800000 : _GEN_134; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_136 = 5'h19 == _T_16[4:0] ? 32'hbe92d7dc : _GEN_135; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_142 = 5'h4 == _T_16[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_143 = 5'h5 == _T_16[4:0] ? 32'hbee5c900 : _GEN_142; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_144 = 5'h6 == _T_16[4:0] ? 32'h80800000 : _GEN_143; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_145 = 5'h7 == _T_16[4:0] ? 32'hbee5c900 : _GEN_144; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_146 = 5'h8 == _T_16[4:0] ? 32'hbf4d57f2 : _GEN_145; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_147 = 5'h9 == _T_16[4:0] ? 32'h80800000 : _GEN_146; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_148 = 5'ha == _T_16[4:0] ? 32'hbf248dba : _GEN_147; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_149 = 5'hb == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_148; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_150 = 5'hc == _T_16[4:0] ? 32'h80800000 : _GEN_149; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_151 = 5'hd == _T_16[4:0] ? 32'hbf4d57f2 : _GEN_150; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_152 = 5'he == _T_16[4:0] ? 32'hbf753ecc : _GEN_151; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_153 = 5'hf == _T_16[4:0] ? 32'h80800000 : _GEN_152; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_154 = 5'h10 == _T_16[4:0] ? 32'hbf6b1034 : _GEN_153; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_155 = 5'h11 == _T_16[4:0] ? 32'hbf3a3528 : _GEN_154; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_156 = 5'h12 == _T_16[4:0] ? 32'h80800000 : _GEN_155; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_157 = 5'h13 == _T_16[4:0] ? 32'hbf7c1c5c : _GEN_156; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_158 = 5'h14 == _T_16[4:0] ? 32'hbeaf1d40 : _GEN_157; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_159 = 5'h15 == _T_16[4:0] ? 32'h80800000 : _GEN_158; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_160 = 5'h16 == _T_16[4:0] ? 32'hbf7f911e : _GEN_159; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_161 = 5'h17 == _T_16[4:0] ? 32'h3dedc210 : _GEN_160; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_162 = 5'h18 == _T_16[4:0] ? 32'h80800000 : _GEN_161; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_163 = 5'h19 == _T_16[4:0] ? 32'hbf753ecc : _GEN_162; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_166 = 5'h1 == _T_16[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_167 = 5'h2 == _T_16[4:0] ? io_in_2_Im : _GEN_166; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_168 = 5'h3 == _T_16[4:0] ? io_in_3_Im : _GEN_167; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_169 = 5'h4 == _T_16[4:0] ? io_in_4_Im : _GEN_168; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_170 = 5'h5 == _T_16[4:0] ? io_in_5_Im : _GEN_169; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_171 = 5'h6 == _T_16[4:0] ? io_in_6_Im : _GEN_170; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_172 = 5'h7 == _T_16[4:0] ? io_in_7_Im : _GEN_171; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_173 = 5'h8 == _T_16[4:0] ? io_in_8_Im : _GEN_172; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_174 = 5'h9 == _T_16[4:0] ? io_in_9_Im : _GEN_173; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_175 = 5'ha == _T_16[4:0] ? io_in_10_Im : _GEN_174; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_176 = 5'hb == _T_16[4:0] ? io_in_11_Im : _GEN_175; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_177 = 5'hc == _T_16[4:0] ? io_in_12_Im : _GEN_176; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_178 = 5'hd == _T_16[4:0] ? io_in_13_Im : _GEN_177; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_179 = 5'he == _T_16[4:0] ? io_in_14_Im : _GEN_178; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_180 = 5'hf == _T_16[4:0] ? io_in_15_Im : _GEN_179; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_181 = 5'h10 == _T_16[4:0] ? io_in_16_Im : _GEN_180; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_182 = 5'h11 == _T_16[4:0] ? io_in_17_Im : _GEN_181; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_183 = 5'h12 == _T_16[4:0] ? io_in_18_Im : _GEN_182; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_184 = 5'h13 == _T_16[4:0] ? io_in_19_Im : _GEN_183; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_185 = 5'h14 == _T_16[4:0] ? io_in_20_Im : _GEN_184; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_186 = 5'h15 == _T_16[4:0] ? io_in_21_Im : _GEN_185; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_187 = 5'h16 == _T_16[4:0] ? io_in_22_Im : _GEN_186; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_188 = 5'h17 == _T_16[4:0] ? io_in_23_Im : _GEN_187; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_189 = 5'h18 == _T_16[4:0] ? io_in_24_Im : _GEN_188; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_190 = 5'h19 == _T_16[4:0] ? io_in_25_Im : _GEN_189; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_193 = 5'h1 == _T_16[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_194 = 5'h2 == _T_16[4:0] ? io_in_2_Re : _GEN_193; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_195 = 5'h3 == _T_16[4:0] ? io_in_3_Re : _GEN_194; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_196 = 5'h4 == _T_16[4:0] ? io_in_4_Re : _GEN_195; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_197 = 5'h5 == _T_16[4:0] ? io_in_5_Re : _GEN_196; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_198 = 5'h6 == _T_16[4:0] ? io_in_6_Re : _GEN_197; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_199 = 5'h7 == _T_16[4:0] ? io_in_7_Re : _GEN_198; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_200 = 5'h8 == _T_16[4:0] ? io_in_8_Re : _GEN_199; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_201 = 5'h9 == _T_16[4:0] ? io_in_9_Re : _GEN_200; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_202 = 5'ha == _T_16[4:0] ? io_in_10_Re : _GEN_201; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_203 = 5'hb == _T_16[4:0] ? io_in_11_Re : _GEN_202; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_204 = 5'hc == _T_16[4:0] ? io_in_12_Re : _GEN_203; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_205 = 5'hd == _T_16[4:0] ? io_in_13_Re : _GEN_204; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_206 = 5'he == _T_16[4:0] ? io_in_14_Re : _GEN_205; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_207 = 5'hf == _T_16[4:0] ? io_in_15_Re : _GEN_206; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_208 = 5'h10 == _T_16[4:0] ? io_in_16_Re : _GEN_207; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_209 = 5'h11 == _T_16[4:0] ? io_in_17_Re : _GEN_208; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_210 = 5'h12 == _T_16[4:0] ? io_in_18_Re : _GEN_209; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_211 = 5'h13 == _T_16[4:0] ? io_in_19_Re : _GEN_210; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_212 = 5'h14 == _T_16[4:0] ? io_in_20_Re : _GEN_211; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_213 = 5'h15 == _T_16[4:0] ? io_in_21_Re : _GEN_212; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_214 = 5'h16 == _T_16[4:0] ? io_in_22_Re : _GEN_213; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_215 = 5'h17 == _T_16[4:0] ? io_in_23_Re : _GEN_214; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_216 = 5'h18 == _T_16[4:0] ? io_in_24_Re : _GEN_215; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_217 = 5'h19 == _T_16[4:0] ? io_in_25_Re : _GEN_216; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_28 = _T_2 + 37'h2; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_223 = 5'h4 == _T_28[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_224 = 5'h5 == _T_28[4:0] ? 32'h3f64c51a : _GEN_223; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_225 = 5'h6 == _T_28[4:0] ? 32'h3f800000 : _GEN_224; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_226 = 5'h7 == _T_28[4:0] ? 32'h3f64c51a : _GEN_225; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_227 = 5'h8 == _T_28[4:0] ? 32'h3f18df62 : _GEN_226; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_228 = 5'h9 == _T_28[4:0] ? 32'h3f800000 : _GEN_227; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_229 = 5'ha == _T_28[4:0] ? 32'h3f441b7c : _GEN_228; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_230 = 5'hb == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_229; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_231 = 5'hc == _T_28[4:0] ? 32'h3f800000 : _GEN_230; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_232 = 5'hd == _T_28[4:0] ? 32'h3f18df62 : _GEN_231; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_233 = 5'he == _T_28[4:0] ? 32'hbe92d7dc : _GEN_232; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_234 = 5'hf == _T_28[4:0] ? 32'h3f800000 : _GEN_233; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_235 = 5'h10 == _T_28[4:0] ? 32'h3ecacaf4 : _GEN_234; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_236 = 5'h11 == _T_28[4:0] ? 32'hbf2fad88 : _GEN_235; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_237 = 5'h12 == _T_28[4:0] ? 32'h3f800000 : _GEN_236; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_238 = 5'h13 == _T_28[4:0] ? 32'h3e31d0d0 : _GEN_237; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_239 = 5'h14 == _T_28[4:0] ? 32'hbf708fb2 : _GEN_238; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_240 = 5'h15 == _T_28[4:0] ? 32'h3f800000 : _GEN_239; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_241 = 5'h16 == _T_28[4:0] ? 32'hbd6e2940 : _GEN_240; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_242 = 5'h17 == _T_28[4:0] ? 32'hbf7e44de : _GEN_241; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_243 = 5'h18 == _T_28[4:0] ? 32'h3f800000 : _GEN_242; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_244 = 5'h19 == _T_28[4:0] ? 32'hbe92d7dc : _GEN_243; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_250 = 5'h4 == _T_28[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_251 = 5'h5 == _T_28[4:0] ? 32'hbee5c900 : _GEN_250; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_252 = 5'h6 == _T_28[4:0] ? 32'h80800000 : _GEN_251; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_253 = 5'h7 == _T_28[4:0] ? 32'hbee5c900 : _GEN_252; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_254 = 5'h8 == _T_28[4:0] ? 32'hbf4d57f2 : _GEN_253; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_255 = 5'h9 == _T_28[4:0] ? 32'h80800000 : _GEN_254; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_256 = 5'ha == _T_28[4:0] ? 32'hbf248dba : _GEN_255; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_257 = 5'hb == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_256; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_258 = 5'hc == _T_28[4:0] ? 32'h80800000 : _GEN_257; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_259 = 5'hd == _T_28[4:0] ? 32'hbf4d57f2 : _GEN_258; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_260 = 5'he == _T_28[4:0] ? 32'hbf753ecc : _GEN_259; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_261 = 5'hf == _T_28[4:0] ? 32'h80800000 : _GEN_260; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_262 = 5'h10 == _T_28[4:0] ? 32'hbf6b1034 : _GEN_261; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_263 = 5'h11 == _T_28[4:0] ? 32'hbf3a3528 : _GEN_262; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_264 = 5'h12 == _T_28[4:0] ? 32'h80800000 : _GEN_263; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_265 = 5'h13 == _T_28[4:0] ? 32'hbf7c1c5c : _GEN_264; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_266 = 5'h14 == _T_28[4:0] ? 32'hbeaf1d40 : _GEN_265; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_267 = 5'h15 == _T_28[4:0] ? 32'h80800000 : _GEN_266; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_268 = 5'h16 == _T_28[4:0] ? 32'hbf7f911e : _GEN_267; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_269 = 5'h17 == _T_28[4:0] ? 32'h3dedc210 : _GEN_268; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_270 = 5'h18 == _T_28[4:0] ? 32'h80800000 : _GEN_269; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_271 = 5'h19 == _T_28[4:0] ? 32'hbf753ecc : _GEN_270; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_274 = 5'h1 == _T_28[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_275 = 5'h2 == _T_28[4:0] ? io_in_2_Im : _GEN_274; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_276 = 5'h3 == _T_28[4:0] ? io_in_3_Im : _GEN_275; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_277 = 5'h4 == _T_28[4:0] ? io_in_4_Im : _GEN_276; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_278 = 5'h5 == _T_28[4:0] ? io_in_5_Im : _GEN_277; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_279 = 5'h6 == _T_28[4:0] ? io_in_6_Im : _GEN_278; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_280 = 5'h7 == _T_28[4:0] ? io_in_7_Im : _GEN_279; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_281 = 5'h8 == _T_28[4:0] ? io_in_8_Im : _GEN_280; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_282 = 5'h9 == _T_28[4:0] ? io_in_9_Im : _GEN_281; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_283 = 5'ha == _T_28[4:0] ? io_in_10_Im : _GEN_282; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_284 = 5'hb == _T_28[4:0] ? io_in_11_Im : _GEN_283; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_285 = 5'hc == _T_28[4:0] ? io_in_12_Im : _GEN_284; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_286 = 5'hd == _T_28[4:0] ? io_in_13_Im : _GEN_285; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_287 = 5'he == _T_28[4:0] ? io_in_14_Im : _GEN_286; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_288 = 5'hf == _T_28[4:0] ? io_in_15_Im : _GEN_287; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_289 = 5'h10 == _T_28[4:0] ? io_in_16_Im : _GEN_288; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_290 = 5'h11 == _T_28[4:0] ? io_in_17_Im : _GEN_289; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_291 = 5'h12 == _T_28[4:0] ? io_in_18_Im : _GEN_290; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_292 = 5'h13 == _T_28[4:0] ? io_in_19_Im : _GEN_291; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_293 = 5'h14 == _T_28[4:0] ? io_in_20_Im : _GEN_292; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_294 = 5'h15 == _T_28[4:0] ? io_in_21_Im : _GEN_293; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_295 = 5'h16 == _T_28[4:0] ? io_in_22_Im : _GEN_294; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_296 = 5'h17 == _T_28[4:0] ? io_in_23_Im : _GEN_295; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_297 = 5'h18 == _T_28[4:0] ? io_in_24_Im : _GEN_296; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_298 = 5'h19 == _T_28[4:0] ? io_in_25_Im : _GEN_297; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_301 = 5'h1 == _T_28[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_302 = 5'h2 == _T_28[4:0] ? io_in_2_Re : _GEN_301; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_303 = 5'h3 == _T_28[4:0] ? io_in_3_Re : _GEN_302; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_304 = 5'h4 == _T_28[4:0] ? io_in_4_Re : _GEN_303; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_305 = 5'h5 == _T_28[4:0] ? io_in_5_Re : _GEN_304; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_306 = 5'h6 == _T_28[4:0] ? io_in_6_Re : _GEN_305; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_307 = 5'h7 == _T_28[4:0] ? io_in_7_Re : _GEN_306; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_308 = 5'h8 == _T_28[4:0] ? io_in_8_Re : _GEN_307; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_309 = 5'h9 == _T_28[4:0] ? io_in_9_Re : _GEN_308; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_310 = 5'ha == _T_28[4:0] ? io_in_10_Re : _GEN_309; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_311 = 5'hb == _T_28[4:0] ? io_in_11_Re : _GEN_310; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_312 = 5'hc == _T_28[4:0] ? io_in_12_Re : _GEN_311; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_313 = 5'hd == _T_28[4:0] ? io_in_13_Re : _GEN_312; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_314 = 5'he == _T_28[4:0] ? io_in_14_Re : _GEN_313; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_315 = 5'hf == _T_28[4:0] ? io_in_15_Re : _GEN_314; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_316 = 5'h10 == _T_28[4:0] ? io_in_16_Re : _GEN_315; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_317 = 5'h11 == _T_28[4:0] ? io_in_17_Re : _GEN_316; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_318 = 5'h12 == _T_28[4:0] ? io_in_18_Re : _GEN_317; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_319 = 5'h13 == _T_28[4:0] ? io_in_19_Re : _GEN_318; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_320 = 5'h14 == _T_28[4:0] ? io_in_20_Re : _GEN_319; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_321 = 5'h15 == _T_28[4:0] ? io_in_21_Re : _GEN_320; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_322 = 5'h16 == _T_28[4:0] ? io_in_22_Re : _GEN_321; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_323 = 5'h17 == _T_28[4:0] ? io_in_23_Re : _GEN_322; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_324 = 5'h18 == _T_28[4:0] ? io_in_24_Re : _GEN_323; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_325 = 5'h19 == _T_28[4:0] ? io_in_25_Re : _GEN_324; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_40 = _T_2 + 37'h3; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_331 = 5'h4 == _T_40[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_332 = 5'h5 == _T_40[4:0] ? 32'h3f64c51a : _GEN_331; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_333 = 5'h6 == _T_40[4:0] ? 32'h3f800000 : _GEN_332; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_334 = 5'h7 == _T_40[4:0] ? 32'h3f64c51a : _GEN_333; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_335 = 5'h8 == _T_40[4:0] ? 32'h3f18df62 : _GEN_334; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_336 = 5'h9 == _T_40[4:0] ? 32'h3f800000 : _GEN_335; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_337 = 5'ha == _T_40[4:0] ? 32'h3f441b7c : _GEN_336; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_338 = 5'hb == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_337; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_339 = 5'hc == _T_40[4:0] ? 32'h3f800000 : _GEN_338; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_340 = 5'hd == _T_40[4:0] ? 32'h3f18df62 : _GEN_339; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_341 = 5'he == _T_40[4:0] ? 32'hbe92d7dc : _GEN_340; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_342 = 5'hf == _T_40[4:0] ? 32'h3f800000 : _GEN_341; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_343 = 5'h10 == _T_40[4:0] ? 32'h3ecacaf4 : _GEN_342; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_344 = 5'h11 == _T_40[4:0] ? 32'hbf2fad88 : _GEN_343; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_345 = 5'h12 == _T_40[4:0] ? 32'h3f800000 : _GEN_344; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_346 = 5'h13 == _T_40[4:0] ? 32'h3e31d0d0 : _GEN_345; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_347 = 5'h14 == _T_40[4:0] ? 32'hbf708fb2 : _GEN_346; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_348 = 5'h15 == _T_40[4:0] ? 32'h3f800000 : _GEN_347; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_349 = 5'h16 == _T_40[4:0] ? 32'hbd6e2940 : _GEN_348; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_350 = 5'h17 == _T_40[4:0] ? 32'hbf7e44de : _GEN_349; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_351 = 5'h18 == _T_40[4:0] ? 32'h3f800000 : _GEN_350; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_352 = 5'h19 == _T_40[4:0] ? 32'hbe92d7dc : _GEN_351; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_358 = 5'h4 == _T_40[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_359 = 5'h5 == _T_40[4:0] ? 32'hbee5c900 : _GEN_358; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_360 = 5'h6 == _T_40[4:0] ? 32'h80800000 : _GEN_359; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_361 = 5'h7 == _T_40[4:0] ? 32'hbee5c900 : _GEN_360; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_362 = 5'h8 == _T_40[4:0] ? 32'hbf4d57f2 : _GEN_361; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_363 = 5'h9 == _T_40[4:0] ? 32'h80800000 : _GEN_362; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_364 = 5'ha == _T_40[4:0] ? 32'hbf248dba : _GEN_363; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_365 = 5'hb == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_364; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_366 = 5'hc == _T_40[4:0] ? 32'h80800000 : _GEN_365; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_367 = 5'hd == _T_40[4:0] ? 32'hbf4d57f2 : _GEN_366; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_368 = 5'he == _T_40[4:0] ? 32'hbf753ecc : _GEN_367; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_369 = 5'hf == _T_40[4:0] ? 32'h80800000 : _GEN_368; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_370 = 5'h10 == _T_40[4:0] ? 32'hbf6b1034 : _GEN_369; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_371 = 5'h11 == _T_40[4:0] ? 32'hbf3a3528 : _GEN_370; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_372 = 5'h12 == _T_40[4:0] ? 32'h80800000 : _GEN_371; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_373 = 5'h13 == _T_40[4:0] ? 32'hbf7c1c5c : _GEN_372; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_374 = 5'h14 == _T_40[4:0] ? 32'hbeaf1d40 : _GEN_373; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_375 = 5'h15 == _T_40[4:0] ? 32'h80800000 : _GEN_374; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_376 = 5'h16 == _T_40[4:0] ? 32'hbf7f911e : _GEN_375; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_377 = 5'h17 == _T_40[4:0] ? 32'h3dedc210 : _GEN_376; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_378 = 5'h18 == _T_40[4:0] ? 32'h80800000 : _GEN_377; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_379 = 5'h19 == _T_40[4:0] ? 32'hbf753ecc : _GEN_378; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_382 = 5'h1 == _T_40[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_383 = 5'h2 == _T_40[4:0] ? io_in_2_Im : _GEN_382; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_384 = 5'h3 == _T_40[4:0] ? io_in_3_Im : _GEN_383; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_385 = 5'h4 == _T_40[4:0] ? io_in_4_Im : _GEN_384; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_386 = 5'h5 == _T_40[4:0] ? io_in_5_Im : _GEN_385; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_387 = 5'h6 == _T_40[4:0] ? io_in_6_Im : _GEN_386; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_388 = 5'h7 == _T_40[4:0] ? io_in_7_Im : _GEN_387; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_389 = 5'h8 == _T_40[4:0] ? io_in_8_Im : _GEN_388; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_390 = 5'h9 == _T_40[4:0] ? io_in_9_Im : _GEN_389; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_391 = 5'ha == _T_40[4:0] ? io_in_10_Im : _GEN_390; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_392 = 5'hb == _T_40[4:0] ? io_in_11_Im : _GEN_391; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_393 = 5'hc == _T_40[4:0] ? io_in_12_Im : _GEN_392; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_394 = 5'hd == _T_40[4:0] ? io_in_13_Im : _GEN_393; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_395 = 5'he == _T_40[4:0] ? io_in_14_Im : _GEN_394; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_396 = 5'hf == _T_40[4:0] ? io_in_15_Im : _GEN_395; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_397 = 5'h10 == _T_40[4:0] ? io_in_16_Im : _GEN_396; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_398 = 5'h11 == _T_40[4:0] ? io_in_17_Im : _GEN_397; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_399 = 5'h12 == _T_40[4:0] ? io_in_18_Im : _GEN_398; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_400 = 5'h13 == _T_40[4:0] ? io_in_19_Im : _GEN_399; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_401 = 5'h14 == _T_40[4:0] ? io_in_20_Im : _GEN_400; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_402 = 5'h15 == _T_40[4:0] ? io_in_21_Im : _GEN_401; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_403 = 5'h16 == _T_40[4:0] ? io_in_22_Im : _GEN_402; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_404 = 5'h17 == _T_40[4:0] ? io_in_23_Im : _GEN_403; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_405 = 5'h18 == _T_40[4:0] ? io_in_24_Im : _GEN_404; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_406 = 5'h19 == _T_40[4:0] ? io_in_25_Im : _GEN_405; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_409 = 5'h1 == _T_40[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_410 = 5'h2 == _T_40[4:0] ? io_in_2_Re : _GEN_409; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_411 = 5'h3 == _T_40[4:0] ? io_in_3_Re : _GEN_410; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_412 = 5'h4 == _T_40[4:0] ? io_in_4_Re : _GEN_411; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_413 = 5'h5 == _T_40[4:0] ? io_in_5_Re : _GEN_412; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_414 = 5'h6 == _T_40[4:0] ? io_in_6_Re : _GEN_413; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_415 = 5'h7 == _T_40[4:0] ? io_in_7_Re : _GEN_414; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_416 = 5'h8 == _T_40[4:0] ? io_in_8_Re : _GEN_415; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_417 = 5'h9 == _T_40[4:0] ? io_in_9_Re : _GEN_416; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_418 = 5'ha == _T_40[4:0] ? io_in_10_Re : _GEN_417; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_419 = 5'hb == _T_40[4:0] ? io_in_11_Re : _GEN_418; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_420 = 5'hc == _T_40[4:0] ? io_in_12_Re : _GEN_419; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_421 = 5'hd == _T_40[4:0] ? io_in_13_Re : _GEN_420; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_422 = 5'he == _T_40[4:0] ? io_in_14_Re : _GEN_421; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_423 = 5'hf == _T_40[4:0] ? io_in_15_Re : _GEN_422; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_424 = 5'h10 == _T_40[4:0] ? io_in_16_Re : _GEN_423; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_425 = 5'h11 == _T_40[4:0] ? io_in_17_Re : _GEN_424; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_426 = 5'h12 == _T_40[4:0] ? io_in_18_Re : _GEN_425; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_427 = 5'h13 == _T_40[4:0] ? io_in_19_Re : _GEN_426; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_428 = 5'h14 == _T_40[4:0] ? io_in_20_Re : _GEN_427; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_429 = 5'h15 == _T_40[4:0] ? io_in_21_Re : _GEN_428; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_430 = 5'h16 == _T_40[4:0] ? io_in_22_Re : _GEN_429; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_431 = 5'h17 == _T_40[4:0] ? io_in_23_Re : _GEN_430; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_432 = 5'h18 == _T_40[4:0] ? io_in_24_Re : _GEN_431; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_433 = 5'h19 == _T_40[4:0] ? io_in_25_Re : _GEN_432; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_52 = _T_2 + 37'h4; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_439 = 5'h4 == _T_52[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_440 = 5'h5 == _T_52[4:0] ? 32'h3f64c51a : _GEN_439; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_441 = 5'h6 == _T_52[4:0] ? 32'h3f800000 : _GEN_440; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_442 = 5'h7 == _T_52[4:0] ? 32'h3f64c51a : _GEN_441; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_443 = 5'h8 == _T_52[4:0] ? 32'h3f18df62 : _GEN_442; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_444 = 5'h9 == _T_52[4:0] ? 32'h3f800000 : _GEN_443; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_445 = 5'ha == _T_52[4:0] ? 32'h3f441b7c : _GEN_444; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_446 = 5'hb == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_445; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_447 = 5'hc == _T_52[4:0] ? 32'h3f800000 : _GEN_446; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_448 = 5'hd == _T_52[4:0] ? 32'h3f18df62 : _GEN_447; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_449 = 5'he == _T_52[4:0] ? 32'hbe92d7dc : _GEN_448; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_450 = 5'hf == _T_52[4:0] ? 32'h3f800000 : _GEN_449; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_451 = 5'h10 == _T_52[4:0] ? 32'h3ecacaf4 : _GEN_450; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_452 = 5'h11 == _T_52[4:0] ? 32'hbf2fad88 : _GEN_451; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_453 = 5'h12 == _T_52[4:0] ? 32'h3f800000 : _GEN_452; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_454 = 5'h13 == _T_52[4:0] ? 32'h3e31d0d0 : _GEN_453; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_455 = 5'h14 == _T_52[4:0] ? 32'hbf708fb2 : _GEN_454; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_456 = 5'h15 == _T_52[4:0] ? 32'h3f800000 : _GEN_455; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_457 = 5'h16 == _T_52[4:0] ? 32'hbd6e2940 : _GEN_456; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_458 = 5'h17 == _T_52[4:0] ? 32'hbf7e44de : _GEN_457; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_459 = 5'h18 == _T_52[4:0] ? 32'h3f800000 : _GEN_458; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_460 = 5'h19 == _T_52[4:0] ? 32'hbe92d7dc : _GEN_459; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_466 = 5'h4 == _T_52[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_467 = 5'h5 == _T_52[4:0] ? 32'hbee5c900 : _GEN_466; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_468 = 5'h6 == _T_52[4:0] ? 32'h80800000 : _GEN_467; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_469 = 5'h7 == _T_52[4:0] ? 32'hbee5c900 : _GEN_468; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_470 = 5'h8 == _T_52[4:0] ? 32'hbf4d57f2 : _GEN_469; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_471 = 5'h9 == _T_52[4:0] ? 32'h80800000 : _GEN_470; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_472 = 5'ha == _T_52[4:0] ? 32'hbf248dba : _GEN_471; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_473 = 5'hb == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_472; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_474 = 5'hc == _T_52[4:0] ? 32'h80800000 : _GEN_473; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_475 = 5'hd == _T_52[4:0] ? 32'hbf4d57f2 : _GEN_474; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_476 = 5'he == _T_52[4:0] ? 32'hbf753ecc : _GEN_475; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_477 = 5'hf == _T_52[4:0] ? 32'h80800000 : _GEN_476; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_478 = 5'h10 == _T_52[4:0] ? 32'hbf6b1034 : _GEN_477; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_479 = 5'h11 == _T_52[4:0] ? 32'hbf3a3528 : _GEN_478; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_480 = 5'h12 == _T_52[4:0] ? 32'h80800000 : _GEN_479; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_481 = 5'h13 == _T_52[4:0] ? 32'hbf7c1c5c : _GEN_480; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_482 = 5'h14 == _T_52[4:0] ? 32'hbeaf1d40 : _GEN_481; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_483 = 5'h15 == _T_52[4:0] ? 32'h80800000 : _GEN_482; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_484 = 5'h16 == _T_52[4:0] ? 32'hbf7f911e : _GEN_483; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_485 = 5'h17 == _T_52[4:0] ? 32'h3dedc210 : _GEN_484; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_486 = 5'h18 == _T_52[4:0] ? 32'h80800000 : _GEN_485; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_487 = 5'h19 == _T_52[4:0] ? 32'hbf753ecc : _GEN_486; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_490 = 5'h1 == _T_52[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_491 = 5'h2 == _T_52[4:0] ? io_in_2_Im : _GEN_490; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_492 = 5'h3 == _T_52[4:0] ? io_in_3_Im : _GEN_491; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_493 = 5'h4 == _T_52[4:0] ? io_in_4_Im : _GEN_492; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_494 = 5'h5 == _T_52[4:0] ? io_in_5_Im : _GEN_493; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_495 = 5'h6 == _T_52[4:0] ? io_in_6_Im : _GEN_494; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_496 = 5'h7 == _T_52[4:0] ? io_in_7_Im : _GEN_495; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_497 = 5'h8 == _T_52[4:0] ? io_in_8_Im : _GEN_496; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_498 = 5'h9 == _T_52[4:0] ? io_in_9_Im : _GEN_497; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_499 = 5'ha == _T_52[4:0] ? io_in_10_Im : _GEN_498; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_500 = 5'hb == _T_52[4:0] ? io_in_11_Im : _GEN_499; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_501 = 5'hc == _T_52[4:0] ? io_in_12_Im : _GEN_500; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_502 = 5'hd == _T_52[4:0] ? io_in_13_Im : _GEN_501; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_503 = 5'he == _T_52[4:0] ? io_in_14_Im : _GEN_502; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_504 = 5'hf == _T_52[4:0] ? io_in_15_Im : _GEN_503; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_505 = 5'h10 == _T_52[4:0] ? io_in_16_Im : _GEN_504; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_506 = 5'h11 == _T_52[4:0] ? io_in_17_Im : _GEN_505; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_507 = 5'h12 == _T_52[4:0] ? io_in_18_Im : _GEN_506; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_508 = 5'h13 == _T_52[4:0] ? io_in_19_Im : _GEN_507; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_509 = 5'h14 == _T_52[4:0] ? io_in_20_Im : _GEN_508; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_510 = 5'h15 == _T_52[4:0] ? io_in_21_Im : _GEN_509; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_511 = 5'h16 == _T_52[4:0] ? io_in_22_Im : _GEN_510; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_512 = 5'h17 == _T_52[4:0] ? io_in_23_Im : _GEN_511; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_513 = 5'h18 == _T_52[4:0] ? io_in_24_Im : _GEN_512; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_514 = 5'h19 == _T_52[4:0] ? io_in_25_Im : _GEN_513; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_517 = 5'h1 == _T_52[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_518 = 5'h2 == _T_52[4:0] ? io_in_2_Re : _GEN_517; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_519 = 5'h3 == _T_52[4:0] ? io_in_3_Re : _GEN_518; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_520 = 5'h4 == _T_52[4:0] ? io_in_4_Re : _GEN_519; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_521 = 5'h5 == _T_52[4:0] ? io_in_5_Re : _GEN_520; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_522 = 5'h6 == _T_52[4:0] ? io_in_6_Re : _GEN_521; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_523 = 5'h7 == _T_52[4:0] ? io_in_7_Re : _GEN_522; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_524 = 5'h8 == _T_52[4:0] ? io_in_8_Re : _GEN_523; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_525 = 5'h9 == _T_52[4:0] ? io_in_9_Re : _GEN_524; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_526 = 5'ha == _T_52[4:0] ? io_in_10_Re : _GEN_525; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_527 = 5'hb == _T_52[4:0] ? io_in_11_Re : _GEN_526; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_528 = 5'hc == _T_52[4:0] ? io_in_12_Re : _GEN_527; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_529 = 5'hd == _T_52[4:0] ? io_in_13_Re : _GEN_528; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_530 = 5'he == _T_52[4:0] ? io_in_14_Re : _GEN_529; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_531 = 5'hf == _T_52[4:0] ? io_in_15_Re : _GEN_530; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_532 = 5'h10 == _T_52[4:0] ? io_in_16_Re : _GEN_531; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_533 = 5'h11 == _T_52[4:0] ? io_in_17_Re : _GEN_532; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_534 = 5'h12 == _T_52[4:0] ? io_in_18_Re : _GEN_533; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_535 = 5'h13 == _T_52[4:0] ? io_in_19_Re : _GEN_534; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_536 = 5'h14 == _T_52[4:0] ? io_in_20_Re : _GEN_535; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_537 = 5'h15 == _T_52[4:0] ? io_in_21_Re : _GEN_536; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_538 = 5'h16 == _T_52[4:0] ? io_in_22_Re : _GEN_537; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_539 = 5'h17 == _T_52[4:0] ? io_in_23_Re : _GEN_538; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_540 = 5'h18 == _T_52[4:0] ? io_in_24_Re : _GEN_539; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_541 = 5'h19 == _T_52[4:0] ? io_in_25_Re : _GEN_540; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_64 = _T_2 + 37'h5; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_547 = 5'h4 == _T_64[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_548 = 5'h5 == _T_64[4:0] ? 32'h3f64c51a : _GEN_547; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_549 = 5'h6 == _T_64[4:0] ? 32'h3f800000 : _GEN_548; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_550 = 5'h7 == _T_64[4:0] ? 32'h3f64c51a : _GEN_549; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_551 = 5'h8 == _T_64[4:0] ? 32'h3f18df62 : _GEN_550; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_552 = 5'h9 == _T_64[4:0] ? 32'h3f800000 : _GEN_551; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_553 = 5'ha == _T_64[4:0] ? 32'h3f441b7c : _GEN_552; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_554 = 5'hb == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_553; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_555 = 5'hc == _T_64[4:0] ? 32'h3f800000 : _GEN_554; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_556 = 5'hd == _T_64[4:0] ? 32'h3f18df62 : _GEN_555; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_557 = 5'he == _T_64[4:0] ? 32'hbe92d7dc : _GEN_556; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_558 = 5'hf == _T_64[4:0] ? 32'h3f800000 : _GEN_557; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_559 = 5'h10 == _T_64[4:0] ? 32'h3ecacaf4 : _GEN_558; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_560 = 5'h11 == _T_64[4:0] ? 32'hbf2fad88 : _GEN_559; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_561 = 5'h12 == _T_64[4:0] ? 32'h3f800000 : _GEN_560; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_562 = 5'h13 == _T_64[4:0] ? 32'h3e31d0d0 : _GEN_561; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_563 = 5'h14 == _T_64[4:0] ? 32'hbf708fb2 : _GEN_562; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_564 = 5'h15 == _T_64[4:0] ? 32'h3f800000 : _GEN_563; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_565 = 5'h16 == _T_64[4:0] ? 32'hbd6e2940 : _GEN_564; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_566 = 5'h17 == _T_64[4:0] ? 32'hbf7e44de : _GEN_565; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_567 = 5'h18 == _T_64[4:0] ? 32'h3f800000 : _GEN_566; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_568 = 5'h19 == _T_64[4:0] ? 32'hbe92d7dc : _GEN_567; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_574 = 5'h4 == _T_64[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_575 = 5'h5 == _T_64[4:0] ? 32'hbee5c900 : _GEN_574; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_576 = 5'h6 == _T_64[4:0] ? 32'h80800000 : _GEN_575; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_577 = 5'h7 == _T_64[4:0] ? 32'hbee5c900 : _GEN_576; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_578 = 5'h8 == _T_64[4:0] ? 32'hbf4d57f2 : _GEN_577; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_579 = 5'h9 == _T_64[4:0] ? 32'h80800000 : _GEN_578; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_580 = 5'ha == _T_64[4:0] ? 32'hbf248dba : _GEN_579; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_581 = 5'hb == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_580; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_582 = 5'hc == _T_64[4:0] ? 32'h80800000 : _GEN_581; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_583 = 5'hd == _T_64[4:0] ? 32'hbf4d57f2 : _GEN_582; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_584 = 5'he == _T_64[4:0] ? 32'hbf753ecc : _GEN_583; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_585 = 5'hf == _T_64[4:0] ? 32'h80800000 : _GEN_584; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_586 = 5'h10 == _T_64[4:0] ? 32'hbf6b1034 : _GEN_585; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_587 = 5'h11 == _T_64[4:0] ? 32'hbf3a3528 : _GEN_586; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_588 = 5'h12 == _T_64[4:0] ? 32'h80800000 : _GEN_587; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_589 = 5'h13 == _T_64[4:0] ? 32'hbf7c1c5c : _GEN_588; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_590 = 5'h14 == _T_64[4:0] ? 32'hbeaf1d40 : _GEN_589; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_591 = 5'h15 == _T_64[4:0] ? 32'h80800000 : _GEN_590; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_592 = 5'h16 == _T_64[4:0] ? 32'hbf7f911e : _GEN_591; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_593 = 5'h17 == _T_64[4:0] ? 32'h3dedc210 : _GEN_592; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_594 = 5'h18 == _T_64[4:0] ? 32'h80800000 : _GEN_593; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_595 = 5'h19 == _T_64[4:0] ? 32'hbf753ecc : _GEN_594; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_598 = 5'h1 == _T_64[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_599 = 5'h2 == _T_64[4:0] ? io_in_2_Im : _GEN_598; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_600 = 5'h3 == _T_64[4:0] ? io_in_3_Im : _GEN_599; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_601 = 5'h4 == _T_64[4:0] ? io_in_4_Im : _GEN_600; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_602 = 5'h5 == _T_64[4:0] ? io_in_5_Im : _GEN_601; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_603 = 5'h6 == _T_64[4:0] ? io_in_6_Im : _GEN_602; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_604 = 5'h7 == _T_64[4:0] ? io_in_7_Im : _GEN_603; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_605 = 5'h8 == _T_64[4:0] ? io_in_8_Im : _GEN_604; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_606 = 5'h9 == _T_64[4:0] ? io_in_9_Im : _GEN_605; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_607 = 5'ha == _T_64[4:0] ? io_in_10_Im : _GEN_606; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_608 = 5'hb == _T_64[4:0] ? io_in_11_Im : _GEN_607; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_609 = 5'hc == _T_64[4:0] ? io_in_12_Im : _GEN_608; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_610 = 5'hd == _T_64[4:0] ? io_in_13_Im : _GEN_609; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_611 = 5'he == _T_64[4:0] ? io_in_14_Im : _GEN_610; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_612 = 5'hf == _T_64[4:0] ? io_in_15_Im : _GEN_611; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_613 = 5'h10 == _T_64[4:0] ? io_in_16_Im : _GEN_612; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_614 = 5'h11 == _T_64[4:0] ? io_in_17_Im : _GEN_613; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_615 = 5'h12 == _T_64[4:0] ? io_in_18_Im : _GEN_614; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_616 = 5'h13 == _T_64[4:0] ? io_in_19_Im : _GEN_615; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_617 = 5'h14 == _T_64[4:0] ? io_in_20_Im : _GEN_616; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_618 = 5'h15 == _T_64[4:0] ? io_in_21_Im : _GEN_617; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_619 = 5'h16 == _T_64[4:0] ? io_in_22_Im : _GEN_618; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_620 = 5'h17 == _T_64[4:0] ? io_in_23_Im : _GEN_619; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_621 = 5'h18 == _T_64[4:0] ? io_in_24_Im : _GEN_620; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_622 = 5'h19 == _T_64[4:0] ? io_in_25_Im : _GEN_621; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_625 = 5'h1 == _T_64[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_626 = 5'h2 == _T_64[4:0] ? io_in_2_Re : _GEN_625; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_627 = 5'h3 == _T_64[4:0] ? io_in_3_Re : _GEN_626; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_628 = 5'h4 == _T_64[4:0] ? io_in_4_Re : _GEN_627; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_629 = 5'h5 == _T_64[4:0] ? io_in_5_Re : _GEN_628; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_630 = 5'h6 == _T_64[4:0] ? io_in_6_Re : _GEN_629; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_631 = 5'h7 == _T_64[4:0] ? io_in_7_Re : _GEN_630; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_632 = 5'h8 == _T_64[4:0] ? io_in_8_Re : _GEN_631; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_633 = 5'h9 == _T_64[4:0] ? io_in_9_Re : _GEN_632; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_634 = 5'ha == _T_64[4:0] ? io_in_10_Re : _GEN_633; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_635 = 5'hb == _T_64[4:0] ? io_in_11_Re : _GEN_634; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_636 = 5'hc == _T_64[4:0] ? io_in_12_Re : _GEN_635; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_637 = 5'hd == _T_64[4:0] ? io_in_13_Re : _GEN_636; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_638 = 5'he == _T_64[4:0] ? io_in_14_Re : _GEN_637; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_639 = 5'hf == _T_64[4:0] ? io_in_15_Re : _GEN_638; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_640 = 5'h10 == _T_64[4:0] ? io_in_16_Re : _GEN_639; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_641 = 5'h11 == _T_64[4:0] ? io_in_17_Re : _GEN_640; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_642 = 5'h12 == _T_64[4:0] ? io_in_18_Re : _GEN_641; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_643 = 5'h13 == _T_64[4:0] ? io_in_19_Re : _GEN_642; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_644 = 5'h14 == _T_64[4:0] ? io_in_20_Re : _GEN_643; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_645 = 5'h15 == _T_64[4:0] ? io_in_21_Re : _GEN_644; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_646 = 5'h16 == _T_64[4:0] ? io_in_22_Re : _GEN_645; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_647 = 5'h17 == _T_64[4:0] ? io_in_23_Re : _GEN_646; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_648 = 5'h18 == _T_64[4:0] ? io_in_24_Re : _GEN_647; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_649 = 5'h19 == _T_64[4:0] ? io_in_25_Re : _GEN_648; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_76 = _T_2 + 37'h6; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_655 = 5'h4 == _T_76[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_656 = 5'h5 == _T_76[4:0] ? 32'h3f64c51a : _GEN_655; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_657 = 5'h6 == _T_76[4:0] ? 32'h3f800000 : _GEN_656; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_658 = 5'h7 == _T_76[4:0] ? 32'h3f64c51a : _GEN_657; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_659 = 5'h8 == _T_76[4:0] ? 32'h3f18df62 : _GEN_658; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_660 = 5'h9 == _T_76[4:0] ? 32'h3f800000 : _GEN_659; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_661 = 5'ha == _T_76[4:0] ? 32'h3f441b7c : _GEN_660; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_662 = 5'hb == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_661; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_663 = 5'hc == _T_76[4:0] ? 32'h3f800000 : _GEN_662; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_664 = 5'hd == _T_76[4:0] ? 32'h3f18df62 : _GEN_663; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_665 = 5'he == _T_76[4:0] ? 32'hbe92d7dc : _GEN_664; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_666 = 5'hf == _T_76[4:0] ? 32'h3f800000 : _GEN_665; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_667 = 5'h10 == _T_76[4:0] ? 32'h3ecacaf4 : _GEN_666; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_668 = 5'h11 == _T_76[4:0] ? 32'hbf2fad88 : _GEN_667; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_669 = 5'h12 == _T_76[4:0] ? 32'h3f800000 : _GEN_668; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_670 = 5'h13 == _T_76[4:0] ? 32'h3e31d0d0 : _GEN_669; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_671 = 5'h14 == _T_76[4:0] ? 32'hbf708fb2 : _GEN_670; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_672 = 5'h15 == _T_76[4:0] ? 32'h3f800000 : _GEN_671; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_673 = 5'h16 == _T_76[4:0] ? 32'hbd6e2940 : _GEN_672; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_674 = 5'h17 == _T_76[4:0] ? 32'hbf7e44de : _GEN_673; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_675 = 5'h18 == _T_76[4:0] ? 32'h3f800000 : _GEN_674; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_676 = 5'h19 == _T_76[4:0] ? 32'hbe92d7dc : _GEN_675; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_682 = 5'h4 == _T_76[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_683 = 5'h5 == _T_76[4:0] ? 32'hbee5c900 : _GEN_682; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_684 = 5'h6 == _T_76[4:0] ? 32'h80800000 : _GEN_683; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_685 = 5'h7 == _T_76[4:0] ? 32'hbee5c900 : _GEN_684; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_686 = 5'h8 == _T_76[4:0] ? 32'hbf4d57f2 : _GEN_685; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_687 = 5'h9 == _T_76[4:0] ? 32'h80800000 : _GEN_686; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_688 = 5'ha == _T_76[4:0] ? 32'hbf248dba : _GEN_687; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_689 = 5'hb == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_688; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_690 = 5'hc == _T_76[4:0] ? 32'h80800000 : _GEN_689; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_691 = 5'hd == _T_76[4:0] ? 32'hbf4d57f2 : _GEN_690; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_692 = 5'he == _T_76[4:0] ? 32'hbf753ecc : _GEN_691; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_693 = 5'hf == _T_76[4:0] ? 32'h80800000 : _GEN_692; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_694 = 5'h10 == _T_76[4:0] ? 32'hbf6b1034 : _GEN_693; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_695 = 5'h11 == _T_76[4:0] ? 32'hbf3a3528 : _GEN_694; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_696 = 5'h12 == _T_76[4:0] ? 32'h80800000 : _GEN_695; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_697 = 5'h13 == _T_76[4:0] ? 32'hbf7c1c5c : _GEN_696; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_698 = 5'h14 == _T_76[4:0] ? 32'hbeaf1d40 : _GEN_697; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_699 = 5'h15 == _T_76[4:0] ? 32'h80800000 : _GEN_698; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_700 = 5'h16 == _T_76[4:0] ? 32'hbf7f911e : _GEN_699; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_701 = 5'h17 == _T_76[4:0] ? 32'h3dedc210 : _GEN_700; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_702 = 5'h18 == _T_76[4:0] ? 32'h80800000 : _GEN_701; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_703 = 5'h19 == _T_76[4:0] ? 32'hbf753ecc : _GEN_702; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_706 = 5'h1 == _T_76[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_707 = 5'h2 == _T_76[4:0] ? io_in_2_Im : _GEN_706; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_708 = 5'h3 == _T_76[4:0] ? io_in_3_Im : _GEN_707; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_709 = 5'h4 == _T_76[4:0] ? io_in_4_Im : _GEN_708; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_710 = 5'h5 == _T_76[4:0] ? io_in_5_Im : _GEN_709; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_711 = 5'h6 == _T_76[4:0] ? io_in_6_Im : _GEN_710; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_712 = 5'h7 == _T_76[4:0] ? io_in_7_Im : _GEN_711; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_713 = 5'h8 == _T_76[4:0] ? io_in_8_Im : _GEN_712; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_714 = 5'h9 == _T_76[4:0] ? io_in_9_Im : _GEN_713; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_715 = 5'ha == _T_76[4:0] ? io_in_10_Im : _GEN_714; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_716 = 5'hb == _T_76[4:0] ? io_in_11_Im : _GEN_715; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_717 = 5'hc == _T_76[4:0] ? io_in_12_Im : _GEN_716; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_718 = 5'hd == _T_76[4:0] ? io_in_13_Im : _GEN_717; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_719 = 5'he == _T_76[4:0] ? io_in_14_Im : _GEN_718; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_720 = 5'hf == _T_76[4:0] ? io_in_15_Im : _GEN_719; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_721 = 5'h10 == _T_76[4:0] ? io_in_16_Im : _GEN_720; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_722 = 5'h11 == _T_76[4:0] ? io_in_17_Im : _GEN_721; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_723 = 5'h12 == _T_76[4:0] ? io_in_18_Im : _GEN_722; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_724 = 5'h13 == _T_76[4:0] ? io_in_19_Im : _GEN_723; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_725 = 5'h14 == _T_76[4:0] ? io_in_20_Im : _GEN_724; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_726 = 5'h15 == _T_76[4:0] ? io_in_21_Im : _GEN_725; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_727 = 5'h16 == _T_76[4:0] ? io_in_22_Im : _GEN_726; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_728 = 5'h17 == _T_76[4:0] ? io_in_23_Im : _GEN_727; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_729 = 5'h18 == _T_76[4:0] ? io_in_24_Im : _GEN_728; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_730 = 5'h19 == _T_76[4:0] ? io_in_25_Im : _GEN_729; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_733 = 5'h1 == _T_76[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_734 = 5'h2 == _T_76[4:0] ? io_in_2_Re : _GEN_733; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_735 = 5'h3 == _T_76[4:0] ? io_in_3_Re : _GEN_734; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_736 = 5'h4 == _T_76[4:0] ? io_in_4_Re : _GEN_735; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_737 = 5'h5 == _T_76[4:0] ? io_in_5_Re : _GEN_736; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_738 = 5'h6 == _T_76[4:0] ? io_in_6_Re : _GEN_737; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_739 = 5'h7 == _T_76[4:0] ? io_in_7_Re : _GEN_738; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_740 = 5'h8 == _T_76[4:0] ? io_in_8_Re : _GEN_739; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_741 = 5'h9 == _T_76[4:0] ? io_in_9_Re : _GEN_740; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_742 = 5'ha == _T_76[4:0] ? io_in_10_Re : _GEN_741; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_743 = 5'hb == _T_76[4:0] ? io_in_11_Re : _GEN_742; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_744 = 5'hc == _T_76[4:0] ? io_in_12_Re : _GEN_743; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_745 = 5'hd == _T_76[4:0] ? io_in_13_Re : _GEN_744; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_746 = 5'he == _T_76[4:0] ? io_in_14_Re : _GEN_745; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_747 = 5'hf == _T_76[4:0] ? io_in_15_Re : _GEN_746; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_748 = 5'h10 == _T_76[4:0] ? io_in_16_Re : _GEN_747; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_749 = 5'h11 == _T_76[4:0] ? io_in_17_Re : _GEN_748; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_750 = 5'h12 == _T_76[4:0] ? io_in_18_Re : _GEN_749; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_751 = 5'h13 == _T_76[4:0] ? io_in_19_Re : _GEN_750; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_752 = 5'h14 == _T_76[4:0] ? io_in_20_Re : _GEN_751; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_753 = 5'h15 == _T_76[4:0] ? io_in_21_Re : _GEN_752; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_754 = 5'h16 == _T_76[4:0] ? io_in_22_Re : _GEN_753; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_755 = 5'h17 == _T_76[4:0] ? io_in_23_Re : _GEN_754; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_756 = 5'h18 == _T_76[4:0] ? io_in_24_Re : _GEN_755; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_757 = 5'h19 == _T_76[4:0] ? io_in_25_Re : _GEN_756; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_88 = _T_2 + 37'h7; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_763 = 5'h4 == _T_88[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_764 = 5'h5 == _T_88[4:0] ? 32'h3f64c51a : _GEN_763; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_765 = 5'h6 == _T_88[4:0] ? 32'h3f800000 : _GEN_764; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_766 = 5'h7 == _T_88[4:0] ? 32'h3f64c51a : _GEN_765; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_767 = 5'h8 == _T_88[4:0] ? 32'h3f18df62 : _GEN_766; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_768 = 5'h9 == _T_88[4:0] ? 32'h3f800000 : _GEN_767; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_769 = 5'ha == _T_88[4:0] ? 32'h3f441b7c : _GEN_768; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_770 = 5'hb == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_769; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_771 = 5'hc == _T_88[4:0] ? 32'h3f800000 : _GEN_770; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_772 = 5'hd == _T_88[4:0] ? 32'h3f18df62 : _GEN_771; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_773 = 5'he == _T_88[4:0] ? 32'hbe92d7dc : _GEN_772; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_774 = 5'hf == _T_88[4:0] ? 32'h3f800000 : _GEN_773; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_775 = 5'h10 == _T_88[4:0] ? 32'h3ecacaf4 : _GEN_774; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_776 = 5'h11 == _T_88[4:0] ? 32'hbf2fad88 : _GEN_775; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_777 = 5'h12 == _T_88[4:0] ? 32'h3f800000 : _GEN_776; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_778 = 5'h13 == _T_88[4:0] ? 32'h3e31d0d0 : _GEN_777; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_779 = 5'h14 == _T_88[4:0] ? 32'hbf708fb2 : _GEN_778; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_780 = 5'h15 == _T_88[4:0] ? 32'h3f800000 : _GEN_779; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_781 = 5'h16 == _T_88[4:0] ? 32'hbd6e2940 : _GEN_780; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_782 = 5'h17 == _T_88[4:0] ? 32'hbf7e44de : _GEN_781; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_783 = 5'h18 == _T_88[4:0] ? 32'h3f800000 : _GEN_782; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_784 = 5'h19 == _T_88[4:0] ? 32'hbe92d7dc : _GEN_783; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_790 = 5'h4 == _T_88[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_791 = 5'h5 == _T_88[4:0] ? 32'hbee5c900 : _GEN_790; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_792 = 5'h6 == _T_88[4:0] ? 32'h80800000 : _GEN_791; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_793 = 5'h7 == _T_88[4:0] ? 32'hbee5c900 : _GEN_792; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_794 = 5'h8 == _T_88[4:0] ? 32'hbf4d57f2 : _GEN_793; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_795 = 5'h9 == _T_88[4:0] ? 32'h80800000 : _GEN_794; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_796 = 5'ha == _T_88[4:0] ? 32'hbf248dba : _GEN_795; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_797 = 5'hb == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_796; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_798 = 5'hc == _T_88[4:0] ? 32'h80800000 : _GEN_797; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_799 = 5'hd == _T_88[4:0] ? 32'hbf4d57f2 : _GEN_798; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_800 = 5'he == _T_88[4:0] ? 32'hbf753ecc : _GEN_799; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_801 = 5'hf == _T_88[4:0] ? 32'h80800000 : _GEN_800; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_802 = 5'h10 == _T_88[4:0] ? 32'hbf6b1034 : _GEN_801; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_803 = 5'h11 == _T_88[4:0] ? 32'hbf3a3528 : _GEN_802; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_804 = 5'h12 == _T_88[4:0] ? 32'h80800000 : _GEN_803; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_805 = 5'h13 == _T_88[4:0] ? 32'hbf7c1c5c : _GEN_804; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_806 = 5'h14 == _T_88[4:0] ? 32'hbeaf1d40 : _GEN_805; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_807 = 5'h15 == _T_88[4:0] ? 32'h80800000 : _GEN_806; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_808 = 5'h16 == _T_88[4:0] ? 32'hbf7f911e : _GEN_807; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_809 = 5'h17 == _T_88[4:0] ? 32'h3dedc210 : _GEN_808; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_810 = 5'h18 == _T_88[4:0] ? 32'h80800000 : _GEN_809; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_811 = 5'h19 == _T_88[4:0] ? 32'hbf753ecc : _GEN_810; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_814 = 5'h1 == _T_88[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_815 = 5'h2 == _T_88[4:0] ? io_in_2_Im : _GEN_814; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_816 = 5'h3 == _T_88[4:0] ? io_in_3_Im : _GEN_815; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_817 = 5'h4 == _T_88[4:0] ? io_in_4_Im : _GEN_816; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_818 = 5'h5 == _T_88[4:0] ? io_in_5_Im : _GEN_817; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_819 = 5'h6 == _T_88[4:0] ? io_in_6_Im : _GEN_818; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_820 = 5'h7 == _T_88[4:0] ? io_in_7_Im : _GEN_819; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_821 = 5'h8 == _T_88[4:0] ? io_in_8_Im : _GEN_820; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_822 = 5'h9 == _T_88[4:0] ? io_in_9_Im : _GEN_821; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_823 = 5'ha == _T_88[4:0] ? io_in_10_Im : _GEN_822; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_824 = 5'hb == _T_88[4:0] ? io_in_11_Im : _GEN_823; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_825 = 5'hc == _T_88[4:0] ? io_in_12_Im : _GEN_824; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_826 = 5'hd == _T_88[4:0] ? io_in_13_Im : _GEN_825; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_827 = 5'he == _T_88[4:0] ? io_in_14_Im : _GEN_826; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_828 = 5'hf == _T_88[4:0] ? io_in_15_Im : _GEN_827; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_829 = 5'h10 == _T_88[4:0] ? io_in_16_Im : _GEN_828; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_830 = 5'h11 == _T_88[4:0] ? io_in_17_Im : _GEN_829; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_831 = 5'h12 == _T_88[4:0] ? io_in_18_Im : _GEN_830; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_832 = 5'h13 == _T_88[4:0] ? io_in_19_Im : _GEN_831; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_833 = 5'h14 == _T_88[4:0] ? io_in_20_Im : _GEN_832; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_834 = 5'h15 == _T_88[4:0] ? io_in_21_Im : _GEN_833; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_835 = 5'h16 == _T_88[4:0] ? io_in_22_Im : _GEN_834; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_836 = 5'h17 == _T_88[4:0] ? io_in_23_Im : _GEN_835; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_837 = 5'h18 == _T_88[4:0] ? io_in_24_Im : _GEN_836; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_838 = 5'h19 == _T_88[4:0] ? io_in_25_Im : _GEN_837; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_841 = 5'h1 == _T_88[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_842 = 5'h2 == _T_88[4:0] ? io_in_2_Re : _GEN_841; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_843 = 5'h3 == _T_88[4:0] ? io_in_3_Re : _GEN_842; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_844 = 5'h4 == _T_88[4:0] ? io_in_4_Re : _GEN_843; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_845 = 5'h5 == _T_88[4:0] ? io_in_5_Re : _GEN_844; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_846 = 5'h6 == _T_88[4:0] ? io_in_6_Re : _GEN_845; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_847 = 5'h7 == _T_88[4:0] ? io_in_7_Re : _GEN_846; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_848 = 5'h8 == _T_88[4:0] ? io_in_8_Re : _GEN_847; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_849 = 5'h9 == _T_88[4:0] ? io_in_9_Re : _GEN_848; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_850 = 5'ha == _T_88[4:0] ? io_in_10_Re : _GEN_849; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_851 = 5'hb == _T_88[4:0] ? io_in_11_Re : _GEN_850; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_852 = 5'hc == _T_88[4:0] ? io_in_12_Re : _GEN_851; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_853 = 5'hd == _T_88[4:0] ? io_in_13_Re : _GEN_852; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_854 = 5'he == _T_88[4:0] ? io_in_14_Re : _GEN_853; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_855 = 5'hf == _T_88[4:0] ? io_in_15_Re : _GEN_854; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_856 = 5'h10 == _T_88[4:0] ? io_in_16_Re : _GEN_855; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_857 = 5'h11 == _T_88[4:0] ? io_in_17_Re : _GEN_856; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_858 = 5'h12 == _T_88[4:0] ? io_in_18_Re : _GEN_857; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_859 = 5'h13 == _T_88[4:0] ? io_in_19_Re : _GEN_858; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_860 = 5'h14 == _T_88[4:0] ? io_in_20_Re : _GEN_859; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_861 = 5'h15 == _T_88[4:0] ? io_in_21_Re : _GEN_860; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_862 = 5'h16 == _T_88[4:0] ? io_in_22_Re : _GEN_861; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_863 = 5'h17 == _T_88[4:0] ? io_in_23_Re : _GEN_862; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_864 = 5'h18 == _T_88[4:0] ? io_in_24_Re : _GEN_863; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_865 = 5'h19 == _T_88[4:0] ? io_in_25_Re : _GEN_864; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_100 = _T_2 + 37'h8; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_871 = 5'h4 == _T_100[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_872 = 5'h5 == _T_100[4:0] ? 32'h3f64c51a : _GEN_871; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_873 = 5'h6 == _T_100[4:0] ? 32'h3f800000 : _GEN_872; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_874 = 5'h7 == _T_100[4:0] ? 32'h3f64c51a : _GEN_873; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_875 = 5'h8 == _T_100[4:0] ? 32'h3f18df62 : _GEN_874; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_876 = 5'h9 == _T_100[4:0] ? 32'h3f800000 : _GEN_875; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_877 = 5'ha == _T_100[4:0] ? 32'h3f441b7c : _GEN_876; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_878 = 5'hb == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_877; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_879 = 5'hc == _T_100[4:0] ? 32'h3f800000 : _GEN_878; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_880 = 5'hd == _T_100[4:0] ? 32'h3f18df62 : _GEN_879; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_881 = 5'he == _T_100[4:0] ? 32'hbe92d7dc : _GEN_880; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_882 = 5'hf == _T_100[4:0] ? 32'h3f800000 : _GEN_881; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_883 = 5'h10 == _T_100[4:0] ? 32'h3ecacaf4 : _GEN_882; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_884 = 5'h11 == _T_100[4:0] ? 32'hbf2fad88 : _GEN_883; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_885 = 5'h12 == _T_100[4:0] ? 32'h3f800000 : _GEN_884; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_886 = 5'h13 == _T_100[4:0] ? 32'h3e31d0d0 : _GEN_885; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_887 = 5'h14 == _T_100[4:0] ? 32'hbf708fb2 : _GEN_886; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_888 = 5'h15 == _T_100[4:0] ? 32'h3f800000 : _GEN_887; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_889 = 5'h16 == _T_100[4:0] ? 32'hbd6e2940 : _GEN_888; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_890 = 5'h17 == _T_100[4:0] ? 32'hbf7e44de : _GEN_889; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_891 = 5'h18 == _T_100[4:0] ? 32'h3f800000 : _GEN_890; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_892 = 5'h19 == _T_100[4:0] ? 32'hbe92d7dc : _GEN_891; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_898 = 5'h4 == _T_100[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_899 = 5'h5 == _T_100[4:0] ? 32'hbee5c900 : _GEN_898; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_900 = 5'h6 == _T_100[4:0] ? 32'h80800000 : _GEN_899; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_901 = 5'h7 == _T_100[4:0] ? 32'hbee5c900 : _GEN_900; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_902 = 5'h8 == _T_100[4:0] ? 32'hbf4d57f2 : _GEN_901; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_903 = 5'h9 == _T_100[4:0] ? 32'h80800000 : _GEN_902; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_904 = 5'ha == _T_100[4:0] ? 32'hbf248dba : _GEN_903; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_905 = 5'hb == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_904; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_906 = 5'hc == _T_100[4:0] ? 32'h80800000 : _GEN_905; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_907 = 5'hd == _T_100[4:0] ? 32'hbf4d57f2 : _GEN_906; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_908 = 5'he == _T_100[4:0] ? 32'hbf753ecc : _GEN_907; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_909 = 5'hf == _T_100[4:0] ? 32'h80800000 : _GEN_908; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_910 = 5'h10 == _T_100[4:0] ? 32'hbf6b1034 : _GEN_909; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_911 = 5'h11 == _T_100[4:0] ? 32'hbf3a3528 : _GEN_910; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_912 = 5'h12 == _T_100[4:0] ? 32'h80800000 : _GEN_911; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_913 = 5'h13 == _T_100[4:0] ? 32'hbf7c1c5c : _GEN_912; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_914 = 5'h14 == _T_100[4:0] ? 32'hbeaf1d40 : _GEN_913; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_915 = 5'h15 == _T_100[4:0] ? 32'h80800000 : _GEN_914; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_916 = 5'h16 == _T_100[4:0] ? 32'hbf7f911e : _GEN_915; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_917 = 5'h17 == _T_100[4:0] ? 32'h3dedc210 : _GEN_916; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_918 = 5'h18 == _T_100[4:0] ? 32'h80800000 : _GEN_917; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_919 = 5'h19 == _T_100[4:0] ? 32'hbf753ecc : _GEN_918; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_922 = 5'h1 == _T_100[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_923 = 5'h2 == _T_100[4:0] ? io_in_2_Im : _GEN_922; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_924 = 5'h3 == _T_100[4:0] ? io_in_3_Im : _GEN_923; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_925 = 5'h4 == _T_100[4:0] ? io_in_4_Im : _GEN_924; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_926 = 5'h5 == _T_100[4:0] ? io_in_5_Im : _GEN_925; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_927 = 5'h6 == _T_100[4:0] ? io_in_6_Im : _GEN_926; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_928 = 5'h7 == _T_100[4:0] ? io_in_7_Im : _GEN_927; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_929 = 5'h8 == _T_100[4:0] ? io_in_8_Im : _GEN_928; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_930 = 5'h9 == _T_100[4:0] ? io_in_9_Im : _GEN_929; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_931 = 5'ha == _T_100[4:0] ? io_in_10_Im : _GEN_930; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_932 = 5'hb == _T_100[4:0] ? io_in_11_Im : _GEN_931; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_933 = 5'hc == _T_100[4:0] ? io_in_12_Im : _GEN_932; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_934 = 5'hd == _T_100[4:0] ? io_in_13_Im : _GEN_933; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_935 = 5'he == _T_100[4:0] ? io_in_14_Im : _GEN_934; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_936 = 5'hf == _T_100[4:0] ? io_in_15_Im : _GEN_935; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_937 = 5'h10 == _T_100[4:0] ? io_in_16_Im : _GEN_936; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_938 = 5'h11 == _T_100[4:0] ? io_in_17_Im : _GEN_937; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_939 = 5'h12 == _T_100[4:0] ? io_in_18_Im : _GEN_938; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_940 = 5'h13 == _T_100[4:0] ? io_in_19_Im : _GEN_939; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_941 = 5'h14 == _T_100[4:0] ? io_in_20_Im : _GEN_940; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_942 = 5'h15 == _T_100[4:0] ? io_in_21_Im : _GEN_941; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_943 = 5'h16 == _T_100[4:0] ? io_in_22_Im : _GEN_942; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_944 = 5'h17 == _T_100[4:0] ? io_in_23_Im : _GEN_943; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_945 = 5'h18 == _T_100[4:0] ? io_in_24_Im : _GEN_944; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_946 = 5'h19 == _T_100[4:0] ? io_in_25_Im : _GEN_945; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_949 = 5'h1 == _T_100[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_950 = 5'h2 == _T_100[4:0] ? io_in_2_Re : _GEN_949; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_951 = 5'h3 == _T_100[4:0] ? io_in_3_Re : _GEN_950; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_952 = 5'h4 == _T_100[4:0] ? io_in_4_Re : _GEN_951; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_953 = 5'h5 == _T_100[4:0] ? io_in_5_Re : _GEN_952; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_954 = 5'h6 == _T_100[4:0] ? io_in_6_Re : _GEN_953; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_955 = 5'h7 == _T_100[4:0] ? io_in_7_Re : _GEN_954; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_956 = 5'h8 == _T_100[4:0] ? io_in_8_Re : _GEN_955; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_957 = 5'h9 == _T_100[4:0] ? io_in_9_Re : _GEN_956; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_958 = 5'ha == _T_100[4:0] ? io_in_10_Re : _GEN_957; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_959 = 5'hb == _T_100[4:0] ? io_in_11_Re : _GEN_958; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_960 = 5'hc == _T_100[4:0] ? io_in_12_Re : _GEN_959; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_961 = 5'hd == _T_100[4:0] ? io_in_13_Re : _GEN_960; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_962 = 5'he == _T_100[4:0] ? io_in_14_Re : _GEN_961; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_963 = 5'hf == _T_100[4:0] ? io_in_15_Re : _GEN_962; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_964 = 5'h10 == _T_100[4:0] ? io_in_16_Re : _GEN_963; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_965 = 5'h11 == _T_100[4:0] ? io_in_17_Re : _GEN_964; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_966 = 5'h12 == _T_100[4:0] ? io_in_18_Re : _GEN_965; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_967 = 5'h13 == _T_100[4:0] ? io_in_19_Re : _GEN_966; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_968 = 5'h14 == _T_100[4:0] ? io_in_20_Re : _GEN_967; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_969 = 5'h15 == _T_100[4:0] ? io_in_21_Re : _GEN_968; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_970 = 5'h16 == _T_100[4:0] ? io_in_22_Re : _GEN_969; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_971 = 5'h17 == _T_100[4:0] ? io_in_23_Re : _GEN_970; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_972 = 5'h18 == _T_100[4:0] ? io_in_24_Re : _GEN_971; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_973 = 5'h19 == _T_100[4:0] ? io_in_25_Re : _GEN_972; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_112 = _T_2 + 37'h9; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_979 = 5'h4 == _T_112[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_980 = 5'h5 == _T_112[4:0] ? 32'h3f64c51a : _GEN_979; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_981 = 5'h6 == _T_112[4:0] ? 32'h3f800000 : _GEN_980; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_982 = 5'h7 == _T_112[4:0] ? 32'h3f64c51a : _GEN_981; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_983 = 5'h8 == _T_112[4:0] ? 32'h3f18df62 : _GEN_982; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_984 = 5'h9 == _T_112[4:0] ? 32'h3f800000 : _GEN_983; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_985 = 5'ha == _T_112[4:0] ? 32'h3f441b7c : _GEN_984; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_986 = 5'hb == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_985; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_987 = 5'hc == _T_112[4:0] ? 32'h3f800000 : _GEN_986; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_988 = 5'hd == _T_112[4:0] ? 32'h3f18df62 : _GEN_987; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_989 = 5'he == _T_112[4:0] ? 32'hbe92d7dc : _GEN_988; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_990 = 5'hf == _T_112[4:0] ? 32'h3f800000 : _GEN_989; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_991 = 5'h10 == _T_112[4:0] ? 32'h3ecacaf4 : _GEN_990; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_992 = 5'h11 == _T_112[4:0] ? 32'hbf2fad88 : _GEN_991; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_993 = 5'h12 == _T_112[4:0] ? 32'h3f800000 : _GEN_992; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_994 = 5'h13 == _T_112[4:0] ? 32'h3e31d0d0 : _GEN_993; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_995 = 5'h14 == _T_112[4:0] ? 32'hbf708fb2 : _GEN_994; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_996 = 5'h15 == _T_112[4:0] ? 32'h3f800000 : _GEN_995; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_997 = 5'h16 == _T_112[4:0] ? 32'hbd6e2940 : _GEN_996; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_998 = 5'h17 == _T_112[4:0] ? 32'hbf7e44de : _GEN_997; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_999 = 5'h18 == _T_112[4:0] ? 32'h3f800000 : _GEN_998; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1000 = 5'h19 == _T_112[4:0] ? 32'hbe92d7dc : _GEN_999; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1006 = 5'h4 == _T_112[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1007 = 5'h5 == _T_112[4:0] ? 32'hbee5c900 : _GEN_1006; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1008 = 5'h6 == _T_112[4:0] ? 32'h80800000 : _GEN_1007; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1009 = 5'h7 == _T_112[4:0] ? 32'hbee5c900 : _GEN_1008; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1010 = 5'h8 == _T_112[4:0] ? 32'hbf4d57f2 : _GEN_1009; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1011 = 5'h9 == _T_112[4:0] ? 32'h80800000 : _GEN_1010; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1012 = 5'ha == _T_112[4:0] ? 32'hbf248dba : _GEN_1011; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1013 = 5'hb == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1012; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1014 = 5'hc == _T_112[4:0] ? 32'h80800000 : _GEN_1013; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1015 = 5'hd == _T_112[4:0] ? 32'hbf4d57f2 : _GEN_1014; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1016 = 5'he == _T_112[4:0] ? 32'hbf753ecc : _GEN_1015; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1017 = 5'hf == _T_112[4:0] ? 32'h80800000 : _GEN_1016; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1018 = 5'h10 == _T_112[4:0] ? 32'hbf6b1034 : _GEN_1017; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1019 = 5'h11 == _T_112[4:0] ? 32'hbf3a3528 : _GEN_1018; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1020 = 5'h12 == _T_112[4:0] ? 32'h80800000 : _GEN_1019; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1021 = 5'h13 == _T_112[4:0] ? 32'hbf7c1c5c : _GEN_1020; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1022 = 5'h14 == _T_112[4:0] ? 32'hbeaf1d40 : _GEN_1021; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1023 = 5'h15 == _T_112[4:0] ? 32'h80800000 : _GEN_1022; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1024 = 5'h16 == _T_112[4:0] ? 32'hbf7f911e : _GEN_1023; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1025 = 5'h17 == _T_112[4:0] ? 32'h3dedc210 : _GEN_1024; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1026 = 5'h18 == _T_112[4:0] ? 32'h80800000 : _GEN_1025; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1027 = 5'h19 == _T_112[4:0] ? 32'hbf753ecc : _GEN_1026; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1030 = 5'h1 == _T_112[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1031 = 5'h2 == _T_112[4:0] ? io_in_2_Im : _GEN_1030; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1032 = 5'h3 == _T_112[4:0] ? io_in_3_Im : _GEN_1031; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1033 = 5'h4 == _T_112[4:0] ? io_in_4_Im : _GEN_1032; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1034 = 5'h5 == _T_112[4:0] ? io_in_5_Im : _GEN_1033; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1035 = 5'h6 == _T_112[4:0] ? io_in_6_Im : _GEN_1034; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1036 = 5'h7 == _T_112[4:0] ? io_in_7_Im : _GEN_1035; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1037 = 5'h8 == _T_112[4:0] ? io_in_8_Im : _GEN_1036; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1038 = 5'h9 == _T_112[4:0] ? io_in_9_Im : _GEN_1037; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1039 = 5'ha == _T_112[4:0] ? io_in_10_Im : _GEN_1038; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1040 = 5'hb == _T_112[4:0] ? io_in_11_Im : _GEN_1039; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1041 = 5'hc == _T_112[4:0] ? io_in_12_Im : _GEN_1040; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1042 = 5'hd == _T_112[4:0] ? io_in_13_Im : _GEN_1041; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1043 = 5'he == _T_112[4:0] ? io_in_14_Im : _GEN_1042; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1044 = 5'hf == _T_112[4:0] ? io_in_15_Im : _GEN_1043; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1045 = 5'h10 == _T_112[4:0] ? io_in_16_Im : _GEN_1044; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1046 = 5'h11 == _T_112[4:0] ? io_in_17_Im : _GEN_1045; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1047 = 5'h12 == _T_112[4:0] ? io_in_18_Im : _GEN_1046; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1048 = 5'h13 == _T_112[4:0] ? io_in_19_Im : _GEN_1047; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1049 = 5'h14 == _T_112[4:0] ? io_in_20_Im : _GEN_1048; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1050 = 5'h15 == _T_112[4:0] ? io_in_21_Im : _GEN_1049; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1051 = 5'h16 == _T_112[4:0] ? io_in_22_Im : _GEN_1050; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1052 = 5'h17 == _T_112[4:0] ? io_in_23_Im : _GEN_1051; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1053 = 5'h18 == _T_112[4:0] ? io_in_24_Im : _GEN_1052; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1054 = 5'h19 == _T_112[4:0] ? io_in_25_Im : _GEN_1053; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1057 = 5'h1 == _T_112[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1058 = 5'h2 == _T_112[4:0] ? io_in_2_Re : _GEN_1057; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1059 = 5'h3 == _T_112[4:0] ? io_in_3_Re : _GEN_1058; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1060 = 5'h4 == _T_112[4:0] ? io_in_4_Re : _GEN_1059; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1061 = 5'h5 == _T_112[4:0] ? io_in_5_Re : _GEN_1060; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1062 = 5'h6 == _T_112[4:0] ? io_in_6_Re : _GEN_1061; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1063 = 5'h7 == _T_112[4:0] ? io_in_7_Re : _GEN_1062; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1064 = 5'h8 == _T_112[4:0] ? io_in_8_Re : _GEN_1063; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1065 = 5'h9 == _T_112[4:0] ? io_in_9_Re : _GEN_1064; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1066 = 5'ha == _T_112[4:0] ? io_in_10_Re : _GEN_1065; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1067 = 5'hb == _T_112[4:0] ? io_in_11_Re : _GEN_1066; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1068 = 5'hc == _T_112[4:0] ? io_in_12_Re : _GEN_1067; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1069 = 5'hd == _T_112[4:0] ? io_in_13_Re : _GEN_1068; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1070 = 5'he == _T_112[4:0] ? io_in_14_Re : _GEN_1069; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1071 = 5'hf == _T_112[4:0] ? io_in_15_Re : _GEN_1070; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1072 = 5'h10 == _T_112[4:0] ? io_in_16_Re : _GEN_1071; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1073 = 5'h11 == _T_112[4:0] ? io_in_17_Re : _GEN_1072; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1074 = 5'h12 == _T_112[4:0] ? io_in_18_Re : _GEN_1073; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1075 = 5'h13 == _T_112[4:0] ? io_in_19_Re : _GEN_1074; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1076 = 5'h14 == _T_112[4:0] ? io_in_20_Re : _GEN_1075; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1077 = 5'h15 == _T_112[4:0] ? io_in_21_Re : _GEN_1076; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1078 = 5'h16 == _T_112[4:0] ? io_in_22_Re : _GEN_1077; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1079 = 5'h17 == _T_112[4:0] ? io_in_23_Re : _GEN_1078; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1080 = 5'h18 == _T_112[4:0] ? io_in_24_Re : _GEN_1079; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1081 = 5'h19 == _T_112[4:0] ? io_in_25_Re : _GEN_1080; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_124 = _T_2 + 37'ha; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1087 = 5'h4 == _T_124[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1088 = 5'h5 == _T_124[4:0] ? 32'h3f64c51a : _GEN_1087; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1089 = 5'h6 == _T_124[4:0] ? 32'h3f800000 : _GEN_1088; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1090 = 5'h7 == _T_124[4:0] ? 32'h3f64c51a : _GEN_1089; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1091 = 5'h8 == _T_124[4:0] ? 32'h3f18df62 : _GEN_1090; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1092 = 5'h9 == _T_124[4:0] ? 32'h3f800000 : _GEN_1091; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1093 = 5'ha == _T_124[4:0] ? 32'h3f441b7c : _GEN_1092; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1094 = 5'hb == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1093; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1095 = 5'hc == _T_124[4:0] ? 32'h3f800000 : _GEN_1094; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1096 = 5'hd == _T_124[4:0] ? 32'h3f18df62 : _GEN_1095; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1097 = 5'he == _T_124[4:0] ? 32'hbe92d7dc : _GEN_1096; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1098 = 5'hf == _T_124[4:0] ? 32'h3f800000 : _GEN_1097; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1099 = 5'h10 == _T_124[4:0] ? 32'h3ecacaf4 : _GEN_1098; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1100 = 5'h11 == _T_124[4:0] ? 32'hbf2fad88 : _GEN_1099; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1101 = 5'h12 == _T_124[4:0] ? 32'h3f800000 : _GEN_1100; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1102 = 5'h13 == _T_124[4:0] ? 32'h3e31d0d0 : _GEN_1101; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1103 = 5'h14 == _T_124[4:0] ? 32'hbf708fb2 : _GEN_1102; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1104 = 5'h15 == _T_124[4:0] ? 32'h3f800000 : _GEN_1103; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1105 = 5'h16 == _T_124[4:0] ? 32'hbd6e2940 : _GEN_1104; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1106 = 5'h17 == _T_124[4:0] ? 32'hbf7e44de : _GEN_1105; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1107 = 5'h18 == _T_124[4:0] ? 32'h3f800000 : _GEN_1106; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1108 = 5'h19 == _T_124[4:0] ? 32'hbe92d7dc : _GEN_1107; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1114 = 5'h4 == _T_124[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1115 = 5'h5 == _T_124[4:0] ? 32'hbee5c900 : _GEN_1114; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1116 = 5'h6 == _T_124[4:0] ? 32'h80800000 : _GEN_1115; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1117 = 5'h7 == _T_124[4:0] ? 32'hbee5c900 : _GEN_1116; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1118 = 5'h8 == _T_124[4:0] ? 32'hbf4d57f2 : _GEN_1117; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1119 = 5'h9 == _T_124[4:0] ? 32'h80800000 : _GEN_1118; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1120 = 5'ha == _T_124[4:0] ? 32'hbf248dba : _GEN_1119; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1121 = 5'hb == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1120; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1122 = 5'hc == _T_124[4:0] ? 32'h80800000 : _GEN_1121; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1123 = 5'hd == _T_124[4:0] ? 32'hbf4d57f2 : _GEN_1122; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1124 = 5'he == _T_124[4:0] ? 32'hbf753ecc : _GEN_1123; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1125 = 5'hf == _T_124[4:0] ? 32'h80800000 : _GEN_1124; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1126 = 5'h10 == _T_124[4:0] ? 32'hbf6b1034 : _GEN_1125; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1127 = 5'h11 == _T_124[4:0] ? 32'hbf3a3528 : _GEN_1126; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1128 = 5'h12 == _T_124[4:0] ? 32'h80800000 : _GEN_1127; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1129 = 5'h13 == _T_124[4:0] ? 32'hbf7c1c5c : _GEN_1128; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1130 = 5'h14 == _T_124[4:0] ? 32'hbeaf1d40 : _GEN_1129; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1131 = 5'h15 == _T_124[4:0] ? 32'h80800000 : _GEN_1130; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1132 = 5'h16 == _T_124[4:0] ? 32'hbf7f911e : _GEN_1131; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1133 = 5'h17 == _T_124[4:0] ? 32'h3dedc210 : _GEN_1132; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1134 = 5'h18 == _T_124[4:0] ? 32'h80800000 : _GEN_1133; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1135 = 5'h19 == _T_124[4:0] ? 32'hbf753ecc : _GEN_1134; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1138 = 5'h1 == _T_124[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1139 = 5'h2 == _T_124[4:0] ? io_in_2_Im : _GEN_1138; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1140 = 5'h3 == _T_124[4:0] ? io_in_3_Im : _GEN_1139; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1141 = 5'h4 == _T_124[4:0] ? io_in_4_Im : _GEN_1140; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1142 = 5'h5 == _T_124[4:0] ? io_in_5_Im : _GEN_1141; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1143 = 5'h6 == _T_124[4:0] ? io_in_6_Im : _GEN_1142; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1144 = 5'h7 == _T_124[4:0] ? io_in_7_Im : _GEN_1143; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1145 = 5'h8 == _T_124[4:0] ? io_in_8_Im : _GEN_1144; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1146 = 5'h9 == _T_124[4:0] ? io_in_9_Im : _GEN_1145; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1147 = 5'ha == _T_124[4:0] ? io_in_10_Im : _GEN_1146; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1148 = 5'hb == _T_124[4:0] ? io_in_11_Im : _GEN_1147; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1149 = 5'hc == _T_124[4:0] ? io_in_12_Im : _GEN_1148; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1150 = 5'hd == _T_124[4:0] ? io_in_13_Im : _GEN_1149; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1151 = 5'he == _T_124[4:0] ? io_in_14_Im : _GEN_1150; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1152 = 5'hf == _T_124[4:0] ? io_in_15_Im : _GEN_1151; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1153 = 5'h10 == _T_124[4:0] ? io_in_16_Im : _GEN_1152; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1154 = 5'h11 == _T_124[4:0] ? io_in_17_Im : _GEN_1153; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1155 = 5'h12 == _T_124[4:0] ? io_in_18_Im : _GEN_1154; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1156 = 5'h13 == _T_124[4:0] ? io_in_19_Im : _GEN_1155; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1157 = 5'h14 == _T_124[4:0] ? io_in_20_Im : _GEN_1156; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1158 = 5'h15 == _T_124[4:0] ? io_in_21_Im : _GEN_1157; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1159 = 5'h16 == _T_124[4:0] ? io_in_22_Im : _GEN_1158; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1160 = 5'h17 == _T_124[4:0] ? io_in_23_Im : _GEN_1159; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1161 = 5'h18 == _T_124[4:0] ? io_in_24_Im : _GEN_1160; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1162 = 5'h19 == _T_124[4:0] ? io_in_25_Im : _GEN_1161; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1165 = 5'h1 == _T_124[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1166 = 5'h2 == _T_124[4:0] ? io_in_2_Re : _GEN_1165; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1167 = 5'h3 == _T_124[4:0] ? io_in_3_Re : _GEN_1166; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1168 = 5'h4 == _T_124[4:0] ? io_in_4_Re : _GEN_1167; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1169 = 5'h5 == _T_124[4:0] ? io_in_5_Re : _GEN_1168; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1170 = 5'h6 == _T_124[4:0] ? io_in_6_Re : _GEN_1169; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1171 = 5'h7 == _T_124[4:0] ? io_in_7_Re : _GEN_1170; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1172 = 5'h8 == _T_124[4:0] ? io_in_8_Re : _GEN_1171; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1173 = 5'h9 == _T_124[4:0] ? io_in_9_Re : _GEN_1172; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1174 = 5'ha == _T_124[4:0] ? io_in_10_Re : _GEN_1173; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1175 = 5'hb == _T_124[4:0] ? io_in_11_Re : _GEN_1174; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1176 = 5'hc == _T_124[4:0] ? io_in_12_Re : _GEN_1175; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1177 = 5'hd == _T_124[4:0] ? io_in_13_Re : _GEN_1176; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1178 = 5'he == _T_124[4:0] ? io_in_14_Re : _GEN_1177; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1179 = 5'hf == _T_124[4:0] ? io_in_15_Re : _GEN_1178; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1180 = 5'h10 == _T_124[4:0] ? io_in_16_Re : _GEN_1179; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1181 = 5'h11 == _T_124[4:0] ? io_in_17_Re : _GEN_1180; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1182 = 5'h12 == _T_124[4:0] ? io_in_18_Re : _GEN_1181; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1183 = 5'h13 == _T_124[4:0] ? io_in_19_Re : _GEN_1182; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1184 = 5'h14 == _T_124[4:0] ? io_in_20_Re : _GEN_1183; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1185 = 5'h15 == _T_124[4:0] ? io_in_21_Re : _GEN_1184; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1186 = 5'h16 == _T_124[4:0] ? io_in_22_Re : _GEN_1185; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1187 = 5'h17 == _T_124[4:0] ? io_in_23_Re : _GEN_1186; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1188 = 5'h18 == _T_124[4:0] ? io_in_24_Re : _GEN_1187; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1189 = 5'h19 == _T_124[4:0] ? io_in_25_Re : _GEN_1188; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_136 = _T_2 + 37'hb; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1195 = 5'h4 == _T_136[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1196 = 5'h5 == _T_136[4:0] ? 32'h3f64c51a : _GEN_1195; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1197 = 5'h6 == _T_136[4:0] ? 32'h3f800000 : _GEN_1196; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1198 = 5'h7 == _T_136[4:0] ? 32'h3f64c51a : _GEN_1197; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1199 = 5'h8 == _T_136[4:0] ? 32'h3f18df62 : _GEN_1198; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1200 = 5'h9 == _T_136[4:0] ? 32'h3f800000 : _GEN_1199; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1201 = 5'ha == _T_136[4:0] ? 32'h3f441b7c : _GEN_1200; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1202 = 5'hb == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1201; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1203 = 5'hc == _T_136[4:0] ? 32'h3f800000 : _GEN_1202; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1204 = 5'hd == _T_136[4:0] ? 32'h3f18df62 : _GEN_1203; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1205 = 5'he == _T_136[4:0] ? 32'hbe92d7dc : _GEN_1204; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1206 = 5'hf == _T_136[4:0] ? 32'h3f800000 : _GEN_1205; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1207 = 5'h10 == _T_136[4:0] ? 32'h3ecacaf4 : _GEN_1206; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1208 = 5'h11 == _T_136[4:0] ? 32'hbf2fad88 : _GEN_1207; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1209 = 5'h12 == _T_136[4:0] ? 32'h3f800000 : _GEN_1208; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1210 = 5'h13 == _T_136[4:0] ? 32'h3e31d0d0 : _GEN_1209; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1211 = 5'h14 == _T_136[4:0] ? 32'hbf708fb2 : _GEN_1210; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1212 = 5'h15 == _T_136[4:0] ? 32'h3f800000 : _GEN_1211; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1213 = 5'h16 == _T_136[4:0] ? 32'hbd6e2940 : _GEN_1212; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1214 = 5'h17 == _T_136[4:0] ? 32'hbf7e44de : _GEN_1213; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1215 = 5'h18 == _T_136[4:0] ? 32'h3f800000 : _GEN_1214; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1216 = 5'h19 == _T_136[4:0] ? 32'hbe92d7dc : _GEN_1215; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1222 = 5'h4 == _T_136[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1223 = 5'h5 == _T_136[4:0] ? 32'hbee5c900 : _GEN_1222; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1224 = 5'h6 == _T_136[4:0] ? 32'h80800000 : _GEN_1223; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1225 = 5'h7 == _T_136[4:0] ? 32'hbee5c900 : _GEN_1224; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1226 = 5'h8 == _T_136[4:0] ? 32'hbf4d57f2 : _GEN_1225; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1227 = 5'h9 == _T_136[4:0] ? 32'h80800000 : _GEN_1226; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1228 = 5'ha == _T_136[4:0] ? 32'hbf248dba : _GEN_1227; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1229 = 5'hb == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1228; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1230 = 5'hc == _T_136[4:0] ? 32'h80800000 : _GEN_1229; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1231 = 5'hd == _T_136[4:0] ? 32'hbf4d57f2 : _GEN_1230; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1232 = 5'he == _T_136[4:0] ? 32'hbf753ecc : _GEN_1231; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1233 = 5'hf == _T_136[4:0] ? 32'h80800000 : _GEN_1232; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1234 = 5'h10 == _T_136[4:0] ? 32'hbf6b1034 : _GEN_1233; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1235 = 5'h11 == _T_136[4:0] ? 32'hbf3a3528 : _GEN_1234; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1236 = 5'h12 == _T_136[4:0] ? 32'h80800000 : _GEN_1235; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1237 = 5'h13 == _T_136[4:0] ? 32'hbf7c1c5c : _GEN_1236; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1238 = 5'h14 == _T_136[4:0] ? 32'hbeaf1d40 : _GEN_1237; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1239 = 5'h15 == _T_136[4:0] ? 32'h80800000 : _GEN_1238; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1240 = 5'h16 == _T_136[4:0] ? 32'hbf7f911e : _GEN_1239; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1241 = 5'h17 == _T_136[4:0] ? 32'h3dedc210 : _GEN_1240; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1242 = 5'h18 == _T_136[4:0] ? 32'h80800000 : _GEN_1241; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1243 = 5'h19 == _T_136[4:0] ? 32'hbf753ecc : _GEN_1242; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1246 = 5'h1 == _T_136[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1247 = 5'h2 == _T_136[4:0] ? io_in_2_Im : _GEN_1246; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1248 = 5'h3 == _T_136[4:0] ? io_in_3_Im : _GEN_1247; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1249 = 5'h4 == _T_136[4:0] ? io_in_4_Im : _GEN_1248; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1250 = 5'h5 == _T_136[4:0] ? io_in_5_Im : _GEN_1249; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1251 = 5'h6 == _T_136[4:0] ? io_in_6_Im : _GEN_1250; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1252 = 5'h7 == _T_136[4:0] ? io_in_7_Im : _GEN_1251; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1253 = 5'h8 == _T_136[4:0] ? io_in_8_Im : _GEN_1252; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1254 = 5'h9 == _T_136[4:0] ? io_in_9_Im : _GEN_1253; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1255 = 5'ha == _T_136[4:0] ? io_in_10_Im : _GEN_1254; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1256 = 5'hb == _T_136[4:0] ? io_in_11_Im : _GEN_1255; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1257 = 5'hc == _T_136[4:0] ? io_in_12_Im : _GEN_1256; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1258 = 5'hd == _T_136[4:0] ? io_in_13_Im : _GEN_1257; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1259 = 5'he == _T_136[4:0] ? io_in_14_Im : _GEN_1258; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1260 = 5'hf == _T_136[4:0] ? io_in_15_Im : _GEN_1259; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1261 = 5'h10 == _T_136[4:0] ? io_in_16_Im : _GEN_1260; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1262 = 5'h11 == _T_136[4:0] ? io_in_17_Im : _GEN_1261; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1263 = 5'h12 == _T_136[4:0] ? io_in_18_Im : _GEN_1262; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1264 = 5'h13 == _T_136[4:0] ? io_in_19_Im : _GEN_1263; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1265 = 5'h14 == _T_136[4:0] ? io_in_20_Im : _GEN_1264; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1266 = 5'h15 == _T_136[4:0] ? io_in_21_Im : _GEN_1265; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1267 = 5'h16 == _T_136[4:0] ? io_in_22_Im : _GEN_1266; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1268 = 5'h17 == _T_136[4:0] ? io_in_23_Im : _GEN_1267; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1269 = 5'h18 == _T_136[4:0] ? io_in_24_Im : _GEN_1268; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1270 = 5'h19 == _T_136[4:0] ? io_in_25_Im : _GEN_1269; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1273 = 5'h1 == _T_136[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1274 = 5'h2 == _T_136[4:0] ? io_in_2_Re : _GEN_1273; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1275 = 5'h3 == _T_136[4:0] ? io_in_3_Re : _GEN_1274; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1276 = 5'h4 == _T_136[4:0] ? io_in_4_Re : _GEN_1275; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1277 = 5'h5 == _T_136[4:0] ? io_in_5_Re : _GEN_1276; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1278 = 5'h6 == _T_136[4:0] ? io_in_6_Re : _GEN_1277; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1279 = 5'h7 == _T_136[4:0] ? io_in_7_Re : _GEN_1278; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1280 = 5'h8 == _T_136[4:0] ? io_in_8_Re : _GEN_1279; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1281 = 5'h9 == _T_136[4:0] ? io_in_9_Re : _GEN_1280; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1282 = 5'ha == _T_136[4:0] ? io_in_10_Re : _GEN_1281; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1283 = 5'hb == _T_136[4:0] ? io_in_11_Re : _GEN_1282; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1284 = 5'hc == _T_136[4:0] ? io_in_12_Re : _GEN_1283; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1285 = 5'hd == _T_136[4:0] ? io_in_13_Re : _GEN_1284; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1286 = 5'he == _T_136[4:0] ? io_in_14_Re : _GEN_1285; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1287 = 5'hf == _T_136[4:0] ? io_in_15_Re : _GEN_1286; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1288 = 5'h10 == _T_136[4:0] ? io_in_16_Re : _GEN_1287; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1289 = 5'h11 == _T_136[4:0] ? io_in_17_Re : _GEN_1288; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1290 = 5'h12 == _T_136[4:0] ? io_in_18_Re : _GEN_1289; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1291 = 5'h13 == _T_136[4:0] ? io_in_19_Re : _GEN_1290; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1292 = 5'h14 == _T_136[4:0] ? io_in_20_Re : _GEN_1291; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1293 = 5'h15 == _T_136[4:0] ? io_in_21_Re : _GEN_1292; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1294 = 5'h16 == _T_136[4:0] ? io_in_22_Re : _GEN_1293; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1295 = 5'h17 == _T_136[4:0] ? io_in_23_Re : _GEN_1294; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1296 = 5'h18 == _T_136[4:0] ? io_in_24_Re : _GEN_1295; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1297 = 5'h19 == _T_136[4:0] ? io_in_25_Re : _GEN_1296; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_148 = _T_2 + 37'hc; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1303 = 5'h4 == _T_148[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1304 = 5'h5 == _T_148[4:0] ? 32'h3f64c51a : _GEN_1303; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1305 = 5'h6 == _T_148[4:0] ? 32'h3f800000 : _GEN_1304; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1306 = 5'h7 == _T_148[4:0] ? 32'h3f64c51a : _GEN_1305; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1307 = 5'h8 == _T_148[4:0] ? 32'h3f18df62 : _GEN_1306; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1308 = 5'h9 == _T_148[4:0] ? 32'h3f800000 : _GEN_1307; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1309 = 5'ha == _T_148[4:0] ? 32'h3f441b7c : _GEN_1308; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1310 = 5'hb == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1309; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1311 = 5'hc == _T_148[4:0] ? 32'h3f800000 : _GEN_1310; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1312 = 5'hd == _T_148[4:0] ? 32'h3f18df62 : _GEN_1311; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1313 = 5'he == _T_148[4:0] ? 32'hbe92d7dc : _GEN_1312; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1314 = 5'hf == _T_148[4:0] ? 32'h3f800000 : _GEN_1313; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1315 = 5'h10 == _T_148[4:0] ? 32'h3ecacaf4 : _GEN_1314; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1316 = 5'h11 == _T_148[4:0] ? 32'hbf2fad88 : _GEN_1315; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1317 = 5'h12 == _T_148[4:0] ? 32'h3f800000 : _GEN_1316; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1318 = 5'h13 == _T_148[4:0] ? 32'h3e31d0d0 : _GEN_1317; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1319 = 5'h14 == _T_148[4:0] ? 32'hbf708fb2 : _GEN_1318; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1320 = 5'h15 == _T_148[4:0] ? 32'h3f800000 : _GEN_1319; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1321 = 5'h16 == _T_148[4:0] ? 32'hbd6e2940 : _GEN_1320; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1322 = 5'h17 == _T_148[4:0] ? 32'hbf7e44de : _GEN_1321; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1323 = 5'h18 == _T_148[4:0] ? 32'h3f800000 : _GEN_1322; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1324 = 5'h19 == _T_148[4:0] ? 32'hbe92d7dc : _GEN_1323; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1330 = 5'h4 == _T_148[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1331 = 5'h5 == _T_148[4:0] ? 32'hbee5c900 : _GEN_1330; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1332 = 5'h6 == _T_148[4:0] ? 32'h80800000 : _GEN_1331; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1333 = 5'h7 == _T_148[4:0] ? 32'hbee5c900 : _GEN_1332; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1334 = 5'h8 == _T_148[4:0] ? 32'hbf4d57f2 : _GEN_1333; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1335 = 5'h9 == _T_148[4:0] ? 32'h80800000 : _GEN_1334; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1336 = 5'ha == _T_148[4:0] ? 32'hbf248dba : _GEN_1335; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1337 = 5'hb == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1336; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1338 = 5'hc == _T_148[4:0] ? 32'h80800000 : _GEN_1337; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1339 = 5'hd == _T_148[4:0] ? 32'hbf4d57f2 : _GEN_1338; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1340 = 5'he == _T_148[4:0] ? 32'hbf753ecc : _GEN_1339; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1341 = 5'hf == _T_148[4:0] ? 32'h80800000 : _GEN_1340; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1342 = 5'h10 == _T_148[4:0] ? 32'hbf6b1034 : _GEN_1341; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1343 = 5'h11 == _T_148[4:0] ? 32'hbf3a3528 : _GEN_1342; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1344 = 5'h12 == _T_148[4:0] ? 32'h80800000 : _GEN_1343; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1345 = 5'h13 == _T_148[4:0] ? 32'hbf7c1c5c : _GEN_1344; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1346 = 5'h14 == _T_148[4:0] ? 32'hbeaf1d40 : _GEN_1345; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1347 = 5'h15 == _T_148[4:0] ? 32'h80800000 : _GEN_1346; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1348 = 5'h16 == _T_148[4:0] ? 32'hbf7f911e : _GEN_1347; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1349 = 5'h17 == _T_148[4:0] ? 32'h3dedc210 : _GEN_1348; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1350 = 5'h18 == _T_148[4:0] ? 32'h80800000 : _GEN_1349; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1351 = 5'h19 == _T_148[4:0] ? 32'hbf753ecc : _GEN_1350; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1354 = 5'h1 == _T_148[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1355 = 5'h2 == _T_148[4:0] ? io_in_2_Im : _GEN_1354; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1356 = 5'h3 == _T_148[4:0] ? io_in_3_Im : _GEN_1355; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1357 = 5'h4 == _T_148[4:0] ? io_in_4_Im : _GEN_1356; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1358 = 5'h5 == _T_148[4:0] ? io_in_5_Im : _GEN_1357; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1359 = 5'h6 == _T_148[4:0] ? io_in_6_Im : _GEN_1358; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1360 = 5'h7 == _T_148[4:0] ? io_in_7_Im : _GEN_1359; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1361 = 5'h8 == _T_148[4:0] ? io_in_8_Im : _GEN_1360; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1362 = 5'h9 == _T_148[4:0] ? io_in_9_Im : _GEN_1361; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1363 = 5'ha == _T_148[4:0] ? io_in_10_Im : _GEN_1362; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1364 = 5'hb == _T_148[4:0] ? io_in_11_Im : _GEN_1363; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1365 = 5'hc == _T_148[4:0] ? io_in_12_Im : _GEN_1364; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1366 = 5'hd == _T_148[4:0] ? io_in_13_Im : _GEN_1365; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1367 = 5'he == _T_148[4:0] ? io_in_14_Im : _GEN_1366; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1368 = 5'hf == _T_148[4:0] ? io_in_15_Im : _GEN_1367; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1369 = 5'h10 == _T_148[4:0] ? io_in_16_Im : _GEN_1368; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1370 = 5'h11 == _T_148[4:0] ? io_in_17_Im : _GEN_1369; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1371 = 5'h12 == _T_148[4:0] ? io_in_18_Im : _GEN_1370; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1372 = 5'h13 == _T_148[4:0] ? io_in_19_Im : _GEN_1371; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1373 = 5'h14 == _T_148[4:0] ? io_in_20_Im : _GEN_1372; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1374 = 5'h15 == _T_148[4:0] ? io_in_21_Im : _GEN_1373; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1375 = 5'h16 == _T_148[4:0] ? io_in_22_Im : _GEN_1374; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1376 = 5'h17 == _T_148[4:0] ? io_in_23_Im : _GEN_1375; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1377 = 5'h18 == _T_148[4:0] ? io_in_24_Im : _GEN_1376; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1378 = 5'h19 == _T_148[4:0] ? io_in_25_Im : _GEN_1377; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1381 = 5'h1 == _T_148[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1382 = 5'h2 == _T_148[4:0] ? io_in_2_Re : _GEN_1381; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1383 = 5'h3 == _T_148[4:0] ? io_in_3_Re : _GEN_1382; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1384 = 5'h4 == _T_148[4:0] ? io_in_4_Re : _GEN_1383; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1385 = 5'h5 == _T_148[4:0] ? io_in_5_Re : _GEN_1384; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1386 = 5'h6 == _T_148[4:0] ? io_in_6_Re : _GEN_1385; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1387 = 5'h7 == _T_148[4:0] ? io_in_7_Re : _GEN_1386; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1388 = 5'h8 == _T_148[4:0] ? io_in_8_Re : _GEN_1387; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1389 = 5'h9 == _T_148[4:0] ? io_in_9_Re : _GEN_1388; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1390 = 5'ha == _T_148[4:0] ? io_in_10_Re : _GEN_1389; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1391 = 5'hb == _T_148[4:0] ? io_in_11_Re : _GEN_1390; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1392 = 5'hc == _T_148[4:0] ? io_in_12_Re : _GEN_1391; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1393 = 5'hd == _T_148[4:0] ? io_in_13_Re : _GEN_1392; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1394 = 5'he == _T_148[4:0] ? io_in_14_Re : _GEN_1393; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1395 = 5'hf == _T_148[4:0] ? io_in_15_Re : _GEN_1394; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1396 = 5'h10 == _T_148[4:0] ? io_in_16_Re : _GEN_1395; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1397 = 5'h11 == _T_148[4:0] ? io_in_17_Re : _GEN_1396; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1398 = 5'h12 == _T_148[4:0] ? io_in_18_Re : _GEN_1397; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1399 = 5'h13 == _T_148[4:0] ? io_in_19_Re : _GEN_1398; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1400 = 5'h14 == _T_148[4:0] ? io_in_20_Re : _GEN_1399; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1401 = 5'h15 == _T_148[4:0] ? io_in_21_Re : _GEN_1400; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1402 = 5'h16 == _T_148[4:0] ? io_in_22_Re : _GEN_1401; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1403 = 5'h17 == _T_148[4:0] ? io_in_23_Re : _GEN_1402; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1404 = 5'h18 == _T_148[4:0] ? io_in_24_Re : _GEN_1403; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1405 = 5'h19 == _T_148[4:0] ? io_in_25_Re : _GEN_1404; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_160 = _T_2 + 37'hd; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1411 = 5'h4 == _T_160[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1412 = 5'h5 == _T_160[4:0] ? 32'h3f64c51a : _GEN_1411; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1413 = 5'h6 == _T_160[4:0] ? 32'h3f800000 : _GEN_1412; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1414 = 5'h7 == _T_160[4:0] ? 32'h3f64c51a : _GEN_1413; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1415 = 5'h8 == _T_160[4:0] ? 32'h3f18df62 : _GEN_1414; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1416 = 5'h9 == _T_160[4:0] ? 32'h3f800000 : _GEN_1415; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1417 = 5'ha == _T_160[4:0] ? 32'h3f441b7c : _GEN_1416; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1418 = 5'hb == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1417; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1419 = 5'hc == _T_160[4:0] ? 32'h3f800000 : _GEN_1418; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1420 = 5'hd == _T_160[4:0] ? 32'h3f18df62 : _GEN_1419; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1421 = 5'he == _T_160[4:0] ? 32'hbe92d7dc : _GEN_1420; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1422 = 5'hf == _T_160[4:0] ? 32'h3f800000 : _GEN_1421; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1423 = 5'h10 == _T_160[4:0] ? 32'h3ecacaf4 : _GEN_1422; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1424 = 5'h11 == _T_160[4:0] ? 32'hbf2fad88 : _GEN_1423; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1425 = 5'h12 == _T_160[4:0] ? 32'h3f800000 : _GEN_1424; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1426 = 5'h13 == _T_160[4:0] ? 32'h3e31d0d0 : _GEN_1425; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1427 = 5'h14 == _T_160[4:0] ? 32'hbf708fb2 : _GEN_1426; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1428 = 5'h15 == _T_160[4:0] ? 32'h3f800000 : _GEN_1427; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1429 = 5'h16 == _T_160[4:0] ? 32'hbd6e2940 : _GEN_1428; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1430 = 5'h17 == _T_160[4:0] ? 32'hbf7e44de : _GEN_1429; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1431 = 5'h18 == _T_160[4:0] ? 32'h3f800000 : _GEN_1430; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1432 = 5'h19 == _T_160[4:0] ? 32'hbe92d7dc : _GEN_1431; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1438 = 5'h4 == _T_160[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1439 = 5'h5 == _T_160[4:0] ? 32'hbee5c900 : _GEN_1438; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1440 = 5'h6 == _T_160[4:0] ? 32'h80800000 : _GEN_1439; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1441 = 5'h7 == _T_160[4:0] ? 32'hbee5c900 : _GEN_1440; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1442 = 5'h8 == _T_160[4:0] ? 32'hbf4d57f2 : _GEN_1441; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1443 = 5'h9 == _T_160[4:0] ? 32'h80800000 : _GEN_1442; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1444 = 5'ha == _T_160[4:0] ? 32'hbf248dba : _GEN_1443; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1445 = 5'hb == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1444; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1446 = 5'hc == _T_160[4:0] ? 32'h80800000 : _GEN_1445; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1447 = 5'hd == _T_160[4:0] ? 32'hbf4d57f2 : _GEN_1446; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1448 = 5'he == _T_160[4:0] ? 32'hbf753ecc : _GEN_1447; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1449 = 5'hf == _T_160[4:0] ? 32'h80800000 : _GEN_1448; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1450 = 5'h10 == _T_160[4:0] ? 32'hbf6b1034 : _GEN_1449; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1451 = 5'h11 == _T_160[4:0] ? 32'hbf3a3528 : _GEN_1450; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1452 = 5'h12 == _T_160[4:0] ? 32'h80800000 : _GEN_1451; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1453 = 5'h13 == _T_160[4:0] ? 32'hbf7c1c5c : _GEN_1452; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1454 = 5'h14 == _T_160[4:0] ? 32'hbeaf1d40 : _GEN_1453; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1455 = 5'h15 == _T_160[4:0] ? 32'h80800000 : _GEN_1454; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1456 = 5'h16 == _T_160[4:0] ? 32'hbf7f911e : _GEN_1455; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1457 = 5'h17 == _T_160[4:0] ? 32'h3dedc210 : _GEN_1456; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1458 = 5'h18 == _T_160[4:0] ? 32'h80800000 : _GEN_1457; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1459 = 5'h19 == _T_160[4:0] ? 32'hbf753ecc : _GEN_1458; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1462 = 5'h1 == _T_160[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1463 = 5'h2 == _T_160[4:0] ? io_in_2_Im : _GEN_1462; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1464 = 5'h3 == _T_160[4:0] ? io_in_3_Im : _GEN_1463; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1465 = 5'h4 == _T_160[4:0] ? io_in_4_Im : _GEN_1464; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1466 = 5'h5 == _T_160[4:0] ? io_in_5_Im : _GEN_1465; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1467 = 5'h6 == _T_160[4:0] ? io_in_6_Im : _GEN_1466; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1468 = 5'h7 == _T_160[4:0] ? io_in_7_Im : _GEN_1467; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1469 = 5'h8 == _T_160[4:0] ? io_in_8_Im : _GEN_1468; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1470 = 5'h9 == _T_160[4:0] ? io_in_9_Im : _GEN_1469; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1471 = 5'ha == _T_160[4:0] ? io_in_10_Im : _GEN_1470; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1472 = 5'hb == _T_160[4:0] ? io_in_11_Im : _GEN_1471; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1473 = 5'hc == _T_160[4:0] ? io_in_12_Im : _GEN_1472; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1474 = 5'hd == _T_160[4:0] ? io_in_13_Im : _GEN_1473; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1475 = 5'he == _T_160[4:0] ? io_in_14_Im : _GEN_1474; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1476 = 5'hf == _T_160[4:0] ? io_in_15_Im : _GEN_1475; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1477 = 5'h10 == _T_160[4:0] ? io_in_16_Im : _GEN_1476; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1478 = 5'h11 == _T_160[4:0] ? io_in_17_Im : _GEN_1477; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1479 = 5'h12 == _T_160[4:0] ? io_in_18_Im : _GEN_1478; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1480 = 5'h13 == _T_160[4:0] ? io_in_19_Im : _GEN_1479; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1481 = 5'h14 == _T_160[4:0] ? io_in_20_Im : _GEN_1480; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1482 = 5'h15 == _T_160[4:0] ? io_in_21_Im : _GEN_1481; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1483 = 5'h16 == _T_160[4:0] ? io_in_22_Im : _GEN_1482; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1484 = 5'h17 == _T_160[4:0] ? io_in_23_Im : _GEN_1483; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1485 = 5'h18 == _T_160[4:0] ? io_in_24_Im : _GEN_1484; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1486 = 5'h19 == _T_160[4:0] ? io_in_25_Im : _GEN_1485; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1489 = 5'h1 == _T_160[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1490 = 5'h2 == _T_160[4:0] ? io_in_2_Re : _GEN_1489; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1491 = 5'h3 == _T_160[4:0] ? io_in_3_Re : _GEN_1490; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1492 = 5'h4 == _T_160[4:0] ? io_in_4_Re : _GEN_1491; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1493 = 5'h5 == _T_160[4:0] ? io_in_5_Re : _GEN_1492; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1494 = 5'h6 == _T_160[4:0] ? io_in_6_Re : _GEN_1493; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1495 = 5'h7 == _T_160[4:0] ? io_in_7_Re : _GEN_1494; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1496 = 5'h8 == _T_160[4:0] ? io_in_8_Re : _GEN_1495; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1497 = 5'h9 == _T_160[4:0] ? io_in_9_Re : _GEN_1496; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1498 = 5'ha == _T_160[4:0] ? io_in_10_Re : _GEN_1497; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1499 = 5'hb == _T_160[4:0] ? io_in_11_Re : _GEN_1498; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1500 = 5'hc == _T_160[4:0] ? io_in_12_Re : _GEN_1499; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1501 = 5'hd == _T_160[4:0] ? io_in_13_Re : _GEN_1500; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1502 = 5'he == _T_160[4:0] ? io_in_14_Re : _GEN_1501; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1503 = 5'hf == _T_160[4:0] ? io_in_15_Re : _GEN_1502; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1504 = 5'h10 == _T_160[4:0] ? io_in_16_Re : _GEN_1503; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1505 = 5'h11 == _T_160[4:0] ? io_in_17_Re : _GEN_1504; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1506 = 5'h12 == _T_160[4:0] ? io_in_18_Re : _GEN_1505; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1507 = 5'h13 == _T_160[4:0] ? io_in_19_Re : _GEN_1506; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1508 = 5'h14 == _T_160[4:0] ? io_in_20_Re : _GEN_1507; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1509 = 5'h15 == _T_160[4:0] ? io_in_21_Re : _GEN_1508; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1510 = 5'h16 == _T_160[4:0] ? io_in_22_Re : _GEN_1509; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1511 = 5'h17 == _T_160[4:0] ? io_in_23_Re : _GEN_1510; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1512 = 5'h18 == _T_160[4:0] ? io_in_24_Re : _GEN_1511; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1513 = 5'h19 == _T_160[4:0] ? io_in_25_Re : _GEN_1512; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_172 = _T_2 + 37'he; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1519 = 5'h4 == _T_172[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1520 = 5'h5 == _T_172[4:0] ? 32'h3f64c51a : _GEN_1519; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1521 = 5'h6 == _T_172[4:0] ? 32'h3f800000 : _GEN_1520; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1522 = 5'h7 == _T_172[4:0] ? 32'h3f64c51a : _GEN_1521; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1523 = 5'h8 == _T_172[4:0] ? 32'h3f18df62 : _GEN_1522; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1524 = 5'h9 == _T_172[4:0] ? 32'h3f800000 : _GEN_1523; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1525 = 5'ha == _T_172[4:0] ? 32'h3f441b7c : _GEN_1524; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1526 = 5'hb == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1525; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1527 = 5'hc == _T_172[4:0] ? 32'h3f800000 : _GEN_1526; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1528 = 5'hd == _T_172[4:0] ? 32'h3f18df62 : _GEN_1527; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1529 = 5'he == _T_172[4:0] ? 32'hbe92d7dc : _GEN_1528; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1530 = 5'hf == _T_172[4:0] ? 32'h3f800000 : _GEN_1529; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1531 = 5'h10 == _T_172[4:0] ? 32'h3ecacaf4 : _GEN_1530; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1532 = 5'h11 == _T_172[4:0] ? 32'hbf2fad88 : _GEN_1531; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1533 = 5'h12 == _T_172[4:0] ? 32'h3f800000 : _GEN_1532; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1534 = 5'h13 == _T_172[4:0] ? 32'h3e31d0d0 : _GEN_1533; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1535 = 5'h14 == _T_172[4:0] ? 32'hbf708fb2 : _GEN_1534; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1536 = 5'h15 == _T_172[4:0] ? 32'h3f800000 : _GEN_1535; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1537 = 5'h16 == _T_172[4:0] ? 32'hbd6e2940 : _GEN_1536; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1538 = 5'h17 == _T_172[4:0] ? 32'hbf7e44de : _GEN_1537; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1539 = 5'h18 == _T_172[4:0] ? 32'h3f800000 : _GEN_1538; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1540 = 5'h19 == _T_172[4:0] ? 32'hbe92d7dc : _GEN_1539; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1546 = 5'h4 == _T_172[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1547 = 5'h5 == _T_172[4:0] ? 32'hbee5c900 : _GEN_1546; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1548 = 5'h6 == _T_172[4:0] ? 32'h80800000 : _GEN_1547; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1549 = 5'h7 == _T_172[4:0] ? 32'hbee5c900 : _GEN_1548; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1550 = 5'h8 == _T_172[4:0] ? 32'hbf4d57f2 : _GEN_1549; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1551 = 5'h9 == _T_172[4:0] ? 32'h80800000 : _GEN_1550; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1552 = 5'ha == _T_172[4:0] ? 32'hbf248dba : _GEN_1551; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1553 = 5'hb == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1552; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1554 = 5'hc == _T_172[4:0] ? 32'h80800000 : _GEN_1553; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1555 = 5'hd == _T_172[4:0] ? 32'hbf4d57f2 : _GEN_1554; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1556 = 5'he == _T_172[4:0] ? 32'hbf753ecc : _GEN_1555; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1557 = 5'hf == _T_172[4:0] ? 32'h80800000 : _GEN_1556; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1558 = 5'h10 == _T_172[4:0] ? 32'hbf6b1034 : _GEN_1557; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1559 = 5'h11 == _T_172[4:0] ? 32'hbf3a3528 : _GEN_1558; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1560 = 5'h12 == _T_172[4:0] ? 32'h80800000 : _GEN_1559; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1561 = 5'h13 == _T_172[4:0] ? 32'hbf7c1c5c : _GEN_1560; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1562 = 5'h14 == _T_172[4:0] ? 32'hbeaf1d40 : _GEN_1561; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1563 = 5'h15 == _T_172[4:0] ? 32'h80800000 : _GEN_1562; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1564 = 5'h16 == _T_172[4:0] ? 32'hbf7f911e : _GEN_1563; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1565 = 5'h17 == _T_172[4:0] ? 32'h3dedc210 : _GEN_1564; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1566 = 5'h18 == _T_172[4:0] ? 32'h80800000 : _GEN_1565; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1567 = 5'h19 == _T_172[4:0] ? 32'hbf753ecc : _GEN_1566; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1570 = 5'h1 == _T_172[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1571 = 5'h2 == _T_172[4:0] ? io_in_2_Im : _GEN_1570; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1572 = 5'h3 == _T_172[4:0] ? io_in_3_Im : _GEN_1571; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1573 = 5'h4 == _T_172[4:0] ? io_in_4_Im : _GEN_1572; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1574 = 5'h5 == _T_172[4:0] ? io_in_5_Im : _GEN_1573; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1575 = 5'h6 == _T_172[4:0] ? io_in_6_Im : _GEN_1574; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1576 = 5'h7 == _T_172[4:0] ? io_in_7_Im : _GEN_1575; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1577 = 5'h8 == _T_172[4:0] ? io_in_8_Im : _GEN_1576; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1578 = 5'h9 == _T_172[4:0] ? io_in_9_Im : _GEN_1577; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1579 = 5'ha == _T_172[4:0] ? io_in_10_Im : _GEN_1578; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1580 = 5'hb == _T_172[4:0] ? io_in_11_Im : _GEN_1579; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1581 = 5'hc == _T_172[4:0] ? io_in_12_Im : _GEN_1580; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1582 = 5'hd == _T_172[4:0] ? io_in_13_Im : _GEN_1581; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1583 = 5'he == _T_172[4:0] ? io_in_14_Im : _GEN_1582; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1584 = 5'hf == _T_172[4:0] ? io_in_15_Im : _GEN_1583; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1585 = 5'h10 == _T_172[4:0] ? io_in_16_Im : _GEN_1584; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1586 = 5'h11 == _T_172[4:0] ? io_in_17_Im : _GEN_1585; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1587 = 5'h12 == _T_172[4:0] ? io_in_18_Im : _GEN_1586; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1588 = 5'h13 == _T_172[4:0] ? io_in_19_Im : _GEN_1587; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1589 = 5'h14 == _T_172[4:0] ? io_in_20_Im : _GEN_1588; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1590 = 5'h15 == _T_172[4:0] ? io_in_21_Im : _GEN_1589; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1591 = 5'h16 == _T_172[4:0] ? io_in_22_Im : _GEN_1590; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1592 = 5'h17 == _T_172[4:0] ? io_in_23_Im : _GEN_1591; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1593 = 5'h18 == _T_172[4:0] ? io_in_24_Im : _GEN_1592; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1594 = 5'h19 == _T_172[4:0] ? io_in_25_Im : _GEN_1593; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1597 = 5'h1 == _T_172[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1598 = 5'h2 == _T_172[4:0] ? io_in_2_Re : _GEN_1597; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1599 = 5'h3 == _T_172[4:0] ? io_in_3_Re : _GEN_1598; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1600 = 5'h4 == _T_172[4:0] ? io_in_4_Re : _GEN_1599; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1601 = 5'h5 == _T_172[4:0] ? io_in_5_Re : _GEN_1600; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1602 = 5'h6 == _T_172[4:0] ? io_in_6_Re : _GEN_1601; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1603 = 5'h7 == _T_172[4:0] ? io_in_7_Re : _GEN_1602; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1604 = 5'h8 == _T_172[4:0] ? io_in_8_Re : _GEN_1603; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1605 = 5'h9 == _T_172[4:0] ? io_in_9_Re : _GEN_1604; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1606 = 5'ha == _T_172[4:0] ? io_in_10_Re : _GEN_1605; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1607 = 5'hb == _T_172[4:0] ? io_in_11_Re : _GEN_1606; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1608 = 5'hc == _T_172[4:0] ? io_in_12_Re : _GEN_1607; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1609 = 5'hd == _T_172[4:0] ? io_in_13_Re : _GEN_1608; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1610 = 5'he == _T_172[4:0] ? io_in_14_Re : _GEN_1609; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1611 = 5'hf == _T_172[4:0] ? io_in_15_Re : _GEN_1610; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1612 = 5'h10 == _T_172[4:0] ? io_in_16_Re : _GEN_1611; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1613 = 5'h11 == _T_172[4:0] ? io_in_17_Re : _GEN_1612; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1614 = 5'h12 == _T_172[4:0] ? io_in_18_Re : _GEN_1613; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1615 = 5'h13 == _T_172[4:0] ? io_in_19_Re : _GEN_1614; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1616 = 5'h14 == _T_172[4:0] ? io_in_20_Re : _GEN_1615; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1617 = 5'h15 == _T_172[4:0] ? io_in_21_Re : _GEN_1616; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1618 = 5'h16 == _T_172[4:0] ? io_in_22_Re : _GEN_1617; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1619 = 5'h17 == _T_172[4:0] ? io_in_23_Re : _GEN_1618; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1620 = 5'h18 == _T_172[4:0] ? io_in_24_Re : _GEN_1619; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1621 = 5'h19 == _T_172[4:0] ? io_in_25_Re : _GEN_1620; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_184 = _T_2 + 37'hf; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1627 = 5'h4 == _T_184[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1628 = 5'h5 == _T_184[4:0] ? 32'h3f64c51a : _GEN_1627; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1629 = 5'h6 == _T_184[4:0] ? 32'h3f800000 : _GEN_1628; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1630 = 5'h7 == _T_184[4:0] ? 32'h3f64c51a : _GEN_1629; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1631 = 5'h8 == _T_184[4:0] ? 32'h3f18df62 : _GEN_1630; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1632 = 5'h9 == _T_184[4:0] ? 32'h3f800000 : _GEN_1631; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1633 = 5'ha == _T_184[4:0] ? 32'h3f441b7c : _GEN_1632; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1634 = 5'hb == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1633; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1635 = 5'hc == _T_184[4:0] ? 32'h3f800000 : _GEN_1634; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1636 = 5'hd == _T_184[4:0] ? 32'h3f18df62 : _GEN_1635; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1637 = 5'he == _T_184[4:0] ? 32'hbe92d7dc : _GEN_1636; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1638 = 5'hf == _T_184[4:0] ? 32'h3f800000 : _GEN_1637; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1639 = 5'h10 == _T_184[4:0] ? 32'h3ecacaf4 : _GEN_1638; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1640 = 5'h11 == _T_184[4:0] ? 32'hbf2fad88 : _GEN_1639; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1641 = 5'h12 == _T_184[4:0] ? 32'h3f800000 : _GEN_1640; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1642 = 5'h13 == _T_184[4:0] ? 32'h3e31d0d0 : _GEN_1641; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1643 = 5'h14 == _T_184[4:0] ? 32'hbf708fb2 : _GEN_1642; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1644 = 5'h15 == _T_184[4:0] ? 32'h3f800000 : _GEN_1643; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1645 = 5'h16 == _T_184[4:0] ? 32'hbd6e2940 : _GEN_1644; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1646 = 5'h17 == _T_184[4:0] ? 32'hbf7e44de : _GEN_1645; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1647 = 5'h18 == _T_184[4:0] ? 32'h3f800000 : _GEN_1646; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1648 = 5'h19 == _T_184[4:0] ? 32'hbe92d7dc : _GEN_1647; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1654 = 5'h4 == _T_184[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1655 = 5'h5 == _T_184[4:0] ? 32'hbee5c900 : _GEN_1654; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1656 = 5'h6 == _T_184[4:0] ? 32'h80800000 : _GEN_1655; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1657 = 5'h7 == _T_184[4:0] ? 32'hbee5c900 : _GEN_1656; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1658 = 5'h8 == _T_184[4:0] ? 32'hbf4d57f2 : _GEN_1657; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1659 = 5'h9 == _T_184[4:0] ? 32'h80800000 : _GEN_1658; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1660 = 5'ha == _T_184[4:0] ? 32'hbf248dba : _GEN_1659; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1661 = 5'hb == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1660; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1662 = 5'hc == _T_184[4:0] ? 32'h80800000 : _GEN_1661; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1663 = 5'hd == _T_184[4:0] ? 32'hbf4d57f2 : _GEN_1662; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1664 = 5'he == _T_184[4:0] ? 32'hbf753ecc : _GEN_1663; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1665 = 5'hf == _T_184[4:0] ? 32'h80800000 : _GEN_1664; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1666 = 5'h10 == _T_184[4:0] ? 32'hbf6b1034 : _GEN_1665; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1667 = 5'h11 == _T_184[4:0] ? 32'hbf3a3528 : _GEN_1666; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1668 = 5'h12 == _T_184[4:0] ? 32'h80800000 : _GEN_1667; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1669 = 5'h13 == _T_184[4:0] ? 32'hbf7c1c5c : _GEN_1668; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1670 = 5'h14 == _T_184[4:0] ? 32'hbeaf1d40 : _GEN_1669; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1671 = 5'h15 == _T_184[4:0] ? 32'h80800000 : _GEN_1670; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1672 = 5'h16 == _T_184[4:0] ? 32'hbf7f911e : _GEN_1671; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1673 = 5'h17 == _T_184[4:0] ? 32'h3dedc210 : _GEN_1672; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1674 = 5'h18 == _T_184[4:0] ? 32'h80800000 : _GEN_1673; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1675 = 5'h19 == _T_184[4:0] ? 32'hbf753ecc : _GEN_1674; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1678 = 5'h1 == _T_184[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1679 = 5'h2 == _T_184[4:0] ? io_in_2_Im : _GEN_1678; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1680 = 5'h3 == _T_184[4:0] ? io_in_3_Im : _GEN_1679; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1681 = 5'h4 == _T_184[4:0] ? io_in_4_Im : _GEN_1680; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1682 = 5'h5 == _T_184[4:0] ? io_in_5_Im : _GEN_1681; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1683 = 5'h6 == _T_184[4:0] ? io_in_6_Im : _GEN_1682; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1684 = 5'h7 == _T_184[4:0] ? io_in_7_Im : _GEN_1683; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1685 = 5'h8 == _T_184[4:0] ? io_in_8_Im : _GEN_1684; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1686 = 5'h9 == _T_184[4:0] ? io_in_9_Im : _GEN_1685; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1687 = 5'ha == _T_184[4:0] ? io_in_10_Im : _GEN_1686; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1688 = 5'hb == _T_184[4:0] ? io_in_11_Im : _GEN_1687; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1689 = 5'hc == _T_184[4:0] ? io_in_12_Im : _GEN_1688; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1690 = 5'hd == _T_184[4:0] ? io_in_13_Im : _GEN_1689; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1691 = 5'he == _T_184[4:0] ? io_in_14_Im : _GEN_1690; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1692 = 5'hf == _T_184[4:0] ? io_in_15_Im : _GEN_1691; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1693 = 5'h10 == _T_184[4:0] ? io_in_16_Im : _GEN_1692; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1694 = 5'h11 == _T_184[4:0] ? io_in_17_Im : _GEN_1693; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1695 = 5'h12 == _T_184[4:0] ? io_in_18_Im : _GEN_1694; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1696 = 5'h13 == _T_184[4:0] ? io_in_19_Im : _GEN_1695; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1697 = 5'h14 == _T_184[4:0] ? io_in_20_Im : _GEN_1696; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1698 = 5'h15 == _T_184[4:0] ? io_in_21_Im : _GEN_1697; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1699 = 5'h16 == _T_184[4:0] ? io_in_22_Im : _GEN_1698; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1700 = 5'h17 == _T_184[4:0] ? io_in_23_Im : _GEN_1699; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1701 = 5'h18 == _T_184[4:0] ? io_in_24_Im : _GEN_1700; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1702 = 5'h19 == _T_184[4:0] ? io_in_25_Im : _GEN_1701; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1705 = 5'h1 == _T_184[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1706 = 5'h2 == _T_184[4:0] ? io_in_2_Re : _GEN_1705; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1707 = 5'h3 == _T_184[4:0] ? io_in_3_Re : _GEN_1706; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1708 = 5'h4 == _T_184[4:0] ? io_in_4_Re : _GEN_1707; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1709 = 5'h5 == _T_184[4:0] ? io_in_5_Re : _GEN_1708; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1710 = 5'h6 == _T_184[4:0] ? io_in_6_Re : _GEN_1709; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1711 = 5'h7 == _T_184[4:0] ? io_in_7_Re : _GEN_1710; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1712 = 5'h8 == _T_184[4:0] ? io_in_8_Re : _GEN_1711; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1713 = 5'h9 == _T_184[4:0] ? io_in_9_Re : _GEN_1712; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1714 = 5'ha == _T_184[4:0] ? io_in_10_Re : _GEN_1713; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1715 = 5'hb == _T_184[4:0] ? io_in_11_Re : _GEN_1714; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1716 = 5'hc == _T_184[4:0] ? io_in_12_Re : _GEN_1715; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1717 = 5'hd == _T_184[4:0] ? io_in_13_Re : _GEN_1716; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1718 = 5'he == _T_184[4:0] ? io_in_14_Re : _GEN_1717; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1719 = 5'hf == _T_184[4:0] ? io_in_15_Re : _GEN_1718; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1720 = 5'h10 == _T_184[4:0] ? io_in_16_Re : _GEN_1719; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1721 = 5'h11 == _T_184[4:0] ? io_in_17_Re : _GEN_1720; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1722 = 5'h12 == _T_184[4:0] ? io_in_18_Re : _GEN_1721; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1723 = 5'h13 == _T_184[4:0] ? io_in_19_Re : _GEN_1722; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1724 = 5'h14 == _T_184[4:0] ? io_in_20_Re : _GEN_1723; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1725 = 5'h15 == _T_184[4:0] ? io_in_21_Re : _GEN_1724; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1726 = 5'h16 == _T_184[4:0] ? io_in_22_Re : _GEN_1725; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1727 = 5'h17 == _T_184[4:0] ? io_in_23_Re : _GEN_1726; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1728 = 5'h18 == _T_184[4:0] ? io_in_24_Re : _GEN_1727; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1729 = 5'h19 == _T_184[4:0] ? io_in_25_Re : _GEN_1728; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_196 = _T_2 + 37'h10; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1735 = 5'h4 == _T_196[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1736 = 5'h5 == _T_196[4:0] ? 32'h3f64c51a : _GEN_1735; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1737 = 5'h6 == _T_196[4:0] ? 32'h3f800000 : _GEN_1736; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1738 = 5'h7 == _T_196[4:0] ? 32'h3f64c51a : _GEN_1737; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1739 = 5'h8 == _T_196[4:0] ? 32'h3f18df62 : _GEN_1738; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1740 = 5'h9 == _T_196[4:0] ? 32'h3f800000 : _GEN_1739; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1741 = 5'ha == _T_196[4:0] ? 32'h3f441b7c : _GEN_1740; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1742 = 5'hb == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1741; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1743 = 5'hc == _T_196[4:0] ? 32'h3f800000 : _GEN_1742; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1744 = 5'hd == _T_196[4:0] ? 32'h3f18df62 : _GEN_1743; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1745 = 5'he == _T_196[4:0] ? 32'hbe92d7dc : _GEN_1744; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1746 = 5'hf == _T_196[4:0] ? 32'h3f800000 : _GEN_1745; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1747 = 5'h10 == _T_196[4:0] ? 32'h3ecacaf4 : _GEN_1746; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1748 = 5'h11 == _T_196[4:0] ? 32'hbf2fad88 : _GEN_1747; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1749 = 5'h12 == _T_196[4:0] ? 32'h3f800000 : _GEN_1748; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1750 = 5'h13 == _T_196[4:0] ? 32'h3e31d0d0 : _GEN_1749; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1751 = 5'h14 == _T_196[4:0] ? 32'hbf708fb2 : _GEN_1750; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1752 = 5'h15 == _T_196[4:0] ? 32'h3f800000 : _GEN_1751; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1753 = 5'h16 == _T_196[4:0] ? 32'hbd6e2940 : _GEN_1752; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1754 = 5'h17 == _T_196[4:0] ? 32'hbf7e44de : _GEN_1753; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1755 = 5'h18 == _T_196[4:0] ? 32'h3f800000 : _GEN_1754; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1756 = 5'h19 == _T_196[4:0] ? 32'hbe92d7dc : _GEN_1755; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1762 = 5'h4 == _T_196[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1763 = 5'h5 == _T_196[4:0] ? 32'hbee5c900 : _GEN_1762; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1764 = 5'h6 == _T_196[4:0] ? 32'h80800000 : _GEN_1763; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1765 = 5'h7 == _T_196[4:0] ? 32'hbee5c900 : _GEN_1764; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1766 = 5'h8 == _T_196[4:0] ? 32'hbf4d57f2 : _GEN_1765; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1767 = 5'h9 == _T_196[4:0] ? 32'h80800000 : _GEN_1766; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1768 = 5'ha == _T_196[4:0] ? 32'hbf248dba : _GEN_1767; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1769 = 5'hb == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1768; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1770 = 5'hc == _T_196[4:0] ? 32'h80800000 : _GEN_1769; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1771 = 5'hd == _T_196[4:0] ? 32'hbf4d57f2 : _GEN_1770; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1772 = 5'he == _T_196[4:0] ? 32'hbf753ecc : _GEN_1771; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1773 = 5'hf == _T_196[4:0] ? 32'h80800000 : _GEN_1772; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1774 = 5'h10 == _T_196[4:0] ? 32'hbf6b1034 : _GEN_1773; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1775 = 5'h11 == _T_196[4:0] ? 32'hbf3a3528 : _GEN_1774; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1776 = 5'h12 == _T_196[4:0] ? 32'h80800000 : _GEN_1775; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1777 = 5'h13 == _T_196[4:0] ? 32'hbf7c1c5c : _GEN_1776; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1778 = 5'h14 == _T_196[4:0] ? 32'hbeaf1d40 : _GEN_1777; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1779 = 5'h15 == _T_196[4:0] ? 32'h80800000 : _GEN_1778; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1780 = 5'h16 == _T_196[4:0] ? 32'hbf7f911e : _GEN_1779; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1781 = 5'h17 == _T_196[4:0] ? 32'h3dedc210 : _GEN_1780; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1782 = 5'h18 == _T_196[4:0] ? 32'h80800000 : _GEN_1781; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1783 = 5'h19 == _T_196[4:0] ? 32'hbf753ecc : _GEN_1782; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1786 = 5'h1 == _T_196[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1787 = 5'h2 == _T_196[4:0] ? io_in_2_Im : _GEN_1786; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1788 = 5'h3 == _T_196[4:0] ? io_in_3_Im : _GEN_1787; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1789 = 5'h4 == _T_196[4:0] ? io_in_4_Im : _GEN_1788; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1790 = 5'h5 == _T_196[4:0] ? io_in_5_Im : _GEN_1789; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1791 = 5'h6 == _T_196[4:0] ? io_in_6_Im : _GEN_1790; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1792 = 5'h7 == _T_196[4:0] ? io_in_7_Im : _GEN_1791; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1793 = 5'h8 == _T_196[4:0] ? io_in_8_Im : _GEN_1792; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1794 = 5'h9 == _T_196[4:0] ? io_in_9_Im : _GEN_1793; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1795 = 5'ha == _T_196[4:0] ? io_in_10_Im : _GEN_1794; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1796 = 5'hb == _T_196[4:0] ? io_in_11_Im : _GEN_1795; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1797 = 5'hc == _T_196[4:0] ? io_in_12_Im : _GEN_1796; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1798 = 5'hd == _T_196[4:0] ? io_in_13_Im : _GEN_1797; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1799 = 5'he == _T_196[4:0] ? io_in_14_Im : _GEN_1798; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1800 = 5'hf == _T_196[4:0] ? io_in_15_Im : _GEN_1799; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1801 = 5'h10 == _T_196[4:0] ? io_in_16_Im : _GEN_1800; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1802 = 5'h11 == _T_196[4:0] ? io_in_17_Im : _GEN_1801; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1803 = 5'h12 == _T_196[4:0] ? io_in_18_Im : _GEN_1802; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1804 = 5'h13 == _T_196[4:0] ? io_in_19_Im : _GEN_1803; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1805 = 5'h14 == _T_196[4:0] ? io_in_20_Im : _GEN_1804; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1806 = 5'h15 == _T_196[4:0] ? io_in_21_Im : _GEN_1805; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1807 = 5'h16 == _T_196[4:0] ? io_in_22_Im : _GEN_1806; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1808 = 5'h17 == _T_196[4:0] ? io_in_23_Im : _GEN_1807; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1809 = 5'h18 == _T_196[4:0] ? io_in_24_Im : _GEN_1808; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1810 = 5'h19 == _T_196[4:0] ? io_in_25_Im : _GEN_1809; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1813 = 5'h1 == _T_196[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1814 = 5'h2 == _T_196[4:0] ? io_in_2_Re : _GEN_1813; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1815 = 5'h3 == _T_196[4:0] ? io_in_3_Re : _GEN_1814; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1816 = 5'h4 == _T_196[4:0] ? io_in_4_Re : _GEN_1815; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1817 = 5'h5 == _T_196[4:0] ? io_in_5_Re : _GEN_1816; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1818 = 5'h6 == _T_196[4:0] ? io_in_6_Re : _GEN_1817; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1819 = 5'h7 == _T_196[4:0] ? io_in_7_Re : _GEN_1818; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1820 = 5'h8 == _T_196[4:0] ? io_in_8_Re : _GEN_1819; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1821 = 5'h9 == _T_196[4:0] ? io_in_9_Re : _GEN_1820; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1822 = 5'ha == _T_196[4:0] ? io_in_10_Re : _GEN_1821; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1823 = 5'hb == _T_196[4:0] ? io_in_11_Re : _GEN_1822; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1824 = 5'hc == _T_196[4:0] ? io_in_12_Re : _GEN_1823; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1825 = 5'hd == _T_196[4:0] ? io_in_13_Re : _GEN_1824; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1826 = 5'he == _T_196[4:0] ? io_in_14_Re : _GEN_1825; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1827 = 5'hf == _T_196[4:0] ? io_in_15_Re : _GEN_1826; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1828 = 5'h10 == _T_196[4:0] ? io_in_16_Re : _GEN_1827; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1829 = 5'h11 == _T_196[4:0] ? io_in_17_Re : _GEN_1828; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1830 = 5'h12 == _T_196[4:0] ? io_in_18_Re : _GEN_1829; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1831 = 5'h13 == _T_196[4:0] ? io_in_19_Re : _GEN_1830; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1832 = 5'h14 == _T_196[4:0] ? io_in_20_Re : _GEN_1831; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1833 = 5'h15 == _T_196[4:0] ? io_in_21_Re : _GEN_1832; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1834 = 5'h16 == _T_196[4:0] ? io_in_22_Re : _GEN_1833; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1835 = 5'h17 == _T_196[4:0] ? io_in_23_Re : _GEN_1834; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1836 = 5'h18 == _T_196[4:0] ? io_in_24_Re : _GEN_1835; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1837 = 5'h19 == _T_196[4:0] ? io_in_25_Re : _GEN_1836; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_208 = _T_2 + 37'h11; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1843 = 5'h4 == _T_208[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1844 = 5'h5 == _T_208[4:0] ? 32'h3f64c51a : _GEN_1843; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1845 = 5'h6 == _T_208[4:0] ? 32'h3f800000 : _GEN_1844; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1846 = 5'h7 == _T_208[4:0] ? 32'h3f64c51a : _GEN_1845; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1847 = 5'h8 == _T_208[4:0] ? 32'h3f18df62 : _GEN_1846; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1848 = 5'h9 == _T_208[4:0] ? 32'h3f800000 : _GEN_1847; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1849 = 5'ha == _T_208[4:0] ? 32'h3f441b7c : _GEN_1848; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1850 = 5'hb == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1849; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1851 = 5'hc == _T_208[4:0] ? 32'h3f800000 : _GEN_1850; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1852 = 5'hd == _T_208[4:0] ? 32'h3f18df62 : _GEN_1851; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1853 = 5'he == _T_208[4:0] ? 32'hbe92d7dc : _GEN_1852; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1854 = 5'hf == _T_208[4:0] ? 32'h3f800000 : _GEN_1853; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1855 = 5'h10 == _T_208[4:0] ? 32'h3ecacaf4 : _GEN_1854; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1856 = 5'h11 == _T_208[4:0] ? 32'hbf2fad88 : _GEN_1855; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1857 = 5'h12 == _T_208[4:0] ? 32'h3f800000 : _GEN_1856; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1858 = 5'h13 == _T_208[4:0] ? 32'h3e31d0d0 : _GEN_1857; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1859 = 5'h14 == _T_208[4:0] ? 32'hbf708fb2 : _GEN_1858; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1860 = 5'h15 == _T_208[4:0] ? 32'h3f800000 : _GEN_1859; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1861 = 5'h16 == _T_208[4:0] ? 32'hbd6e2940 : _GEN_1860; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1862 = 5'h17 == _T_208[4:0] ? 32'hbf7e44de : _GEN_1861; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1863 = 5'h18 == _T_208[4:0] ? 32'h3f800000 : _GEN_1862; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1864 = 5'h19 == _T_208[4:0] ? 32'hbe92d7dc : _GEN_1863; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1870 = 5'h4 == _T_208[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1871 = 5'h5 == _T_208[4:0] ? 32'hbee5c900 : _GEN_1870; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1872 = 5'h6 == _T_208[4:0] ? 32'h80800000 : _GEN_1871; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1873 = 5'h7 == _T_208[4:0] ? 32'hbee5c900 : _GEN_1872; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1874 = 5'h8 == _T_208[4:0] ? 32'hbf4d57f2 : _GEN_1873; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1875 = 5'h9 == _T_208[4:0] ? 32'h80800000 : _GEN_1874; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1876 = 5'ha == _T_208[4:0] ? 32'hbf248dba : _GEN_1875; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1877 = 5'hb == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1876; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1878 = 5'hc == _T_208[4:0] ? 32'h80800000 : _GEN_1877; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1879 = 5'hd == _T_208[4:0] ? 32'hbf4d57f2 : _GEN_1878; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1880 = 5'he == _T_208[4:0] ? 32'hbf753ecc : _GEN_1879; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1881 = 5'hf == _T_208[4:0] ? 32'h80800000 : _GEN_1880; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1882 = 5'h10 == _T_208[4:0] ? 32'hbf6b1034 : _GEN_1881; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1883 = 5'h11 == _T_208[4:0] ? 32'hbf3a3528 : _GEN_1882; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1884 = 5'h12 == _T_208[4:0] ? 32'h80800000 : _GEN_1883; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1885 = 5'h13 == _T_208[4:0] ? 32'hbf7c1c5c : _GEN_1884; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1886 = 5'h14 == _T_208[4:0] ? 32'hbeaf1d40 : _GEN_1885; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1887 = 5'h15 == _T_208[4:0] ? 32'h80800000 : _GEN_1886; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1888 = 5'h16 == _T_208[4:0] ? 32'hbf7f911e : _GEN_1887; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1889 = 5'h17 == _T_208[4:0] ? 32'h3dedc210 : _GEN_1888; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1890 = 5'h18 == _T_208[4:0] ? 32'h80800000 : _GEN_1889; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1891 = 5'h19 == _T_208[4:0] ? 32'hbf753ecc : _GEN_1890; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1894 = 5'h1 == _T_208[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1895 = 5'h2 == _T_208[4:0] ? io_in_2_Im : _GEN_1894; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1896 = 5'h3 == _T_208[4:0] ? io_in_3_Im : _GEN_1895; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1897 = 5'h4 == _T_208[4:0] ? io_in_4_Im : _GEN_1896; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1898 = 5'h5 == _T_208[4:0] ? io_in_5_Im : _GEN_1897; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1899 = 5'h6 == _T_208[4:0] ? io_in_6_Im : _GEN_1898; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1900 = 5'h7 == _T_208[4:0] ? io_in_7_Im : _GEN_1899; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1901 = 5'h8 == _T_208[4:0] ? io_in_8_Im : _GEN_1900; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1902 = 5'h9 == _T_208[4:0] ? io_in_9_Im : _GEN_1901; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1903 = 5'ha == _T_208[4:0] ? io_in_10_Im : _GEN_1902; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1904 = 5'hb == _T_208[4:0] ? io_in_11_Im : _GEN_1903; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1905 = 5'hc == _T_208[4:0] ? io_in_12_Im : _GEN_1904; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1906 = 5'hd == _T_208[4:0] ? io_in_13_Im : _GEN_1905; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1907 = 5'he == _T_208[4:0] ? io_in_14_Im : _GEN_1906; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1908 = 5'hf == _T_208[4:0] ? io_in_15_Im : _GEN_1907; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1909 = 5'h10 == _T_208[4:0] ? io_in_16_Im : _GEN_1908; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1910 = 5'h11 == _T_208[4:0] ? io_in_17_Im : _GEN_1909; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1911 = 5'h12 == _T_208[4:0] ? io_in_18_Im : _GEN_1910; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1912 = 5'h13 == _T_208[4:0] ? io_in_19_Im : _GEN_1911; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1913 = 5'h14 == _T_208[4:0] ? io_in_20_Im : _GEN_1912; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1914 = 5'h15 == _T_208[4:0] ? io_in_21_Im : _GEN_1913; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1915 = 5'h16 == _T_208[4:0] ? io_in_22_Im : _GEN_1914; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1916 = 5'h17 == _T_208[4:0] ? io_in_23_Im : _GEN_1915; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1917 = 5'h18 == _T_208[4:0] ? io_in_24_Im : _GEN_1916; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1918 = 5'h19 == _T_208[4:0] ? io_in_25_Im : _GEN_1917; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1921 = 5'h1 == _T_208[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1922 = 5'h2 == _T_208[4:0] ? io_in_2_Re : _GEN_1921; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1923 = 5'h3 == _T_208[4:0] ? io_in_3_Re : _GEN_1922; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1924 = 5'h4 == _T_208[4:0] ? io_in_4_Re : _GEN_1923; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1925 = 5'h5 == _T_208[4:0] ? io_in_5_Re : _GEN_1924; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1926 = 5'h6 == _T_208[4:0] ? io_in_6_Re : _GEN_1925; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1927 = 5'h7 == _T_208[4:0] ? io_in_7_Re : _GEN_1926; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1928 = 5'h8 == _T_208[4:0] ? io_in_8_Re : _GEN_1927; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1929 = 5'h9 == _T_208[4:0] ? io_in_9_Re : _GEN_1928; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1930 = 5'ha == _T_208[4:0] ? io_in_10_Re : _GEN_1929; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1931 = 5'hb == _T_208[4:0] ? io_in_11_Re : _GEN_1930; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1932 = 5'hc == _T_208[4:0] ? io_in_12_Re : _GEN_1931; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1933 = 5'hd == _T_208[4:0] ? io_in_13_Re : _GEN_1932; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1934 = 5'he == _T_208[4:0] ? io_in_14_Re : _GEN_1933; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1935 = 5'hf == _T_208[4:0] ? io_in_15_Re : _GEN_1934; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1936 = 5'h10 == _T_208[4:0] ? io_in_16_Re : _GEN_1935; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1937 = 5'h11 == _T_208[4:0] ? io_in_17_Re : _GEN_1936; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1938 = 5'h12 == _T_208[4:0] ? io_in_18_Re : _GEN_1937; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1939 = 5'h13 == _T_208[4:0] ? io_in_19_Re : _GEN_1938; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1940 = 5'h14 == _T_208[4:0] ? io_in_20_Re : _GEN_1939; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1941 = 5'h15 == _T_208[4:0] ? io_in_21_Re : _GEN_1940; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1942 = 5'h16 == _T_208[4:0] ? io_in_22_Re : _GEN_1941; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1943 = 5'h17 == _T_208[4:0] ? io_in_23_Re : _GEN_1942; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1944 = 5'h18 == _T_208[4:0] ? io_in_24_Re : _GEN_1943; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_1945 = 5'h19 == _T_208[4:0] ? io_in_25_Re : _GEN_1944; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_220 = _T_2 + 37'h12; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_1951 = 5'h4 == _T_220[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1952 = 5'h5 == _T_220[4:0] ? 32'h3f64c51a : _GEN_1951; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1953 = 5'h6 == _T_220[4:0] ? 32'h3f800000 : _GEN_1952; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1954 = 5'h7 == _T_220[4:0] ? 32'h3f64c51a : _GEN_1953; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1955 = 5'h8 == _T_220[4:0] ? 32'h3f18df62 : _GEN_1954; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1956 = 5'h9 == _T_220[4:0] ? 32'h3f800000 : _GEN_1955; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1957 = 5'ha == _T_220[4:0] ? 32'h3f441b7c : _GEN_1956; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1958 = 5'hb == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1957; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1959 = 5'hc == _T_220[4:0] ? 32'h3f800000 : _GEN_1958; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1960 = 5'hd == _T_220[4:0] ? 32'h3f18df62 : _GEN_1959; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1961 = 5'he == _T_220[4:0] ? 32'hbe92d7dc : _GEN_1960; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1962 = 5'hf == _T_220[4:0] ? 32'h3f800000 : _GEN_1961; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1963 = 5'h10 == _T_220[4:0] ? 32'h3ecacaf4 : _GEN_1962; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1964 = 5'h11 == _T_220[4:0] ? 32'hbf2fad88 : _GEN_1963; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1965 = 5'h12 == _T_220[4:0] ? 32'h3f800000 : _GEN_1964; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1966 = 5'h13 == _T_220[4:0] ? 32'h3e31d0d0 : _GEN_1965; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1967 = 5'h14 == _T_220[4:0] ? 32'hbf708fb2 : _GEN_1966; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1968 = 5'h15 == _T_220[4:0] ? 32'h3f800000 : _GEN_1967; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1969 = 5'h16 == _T_220[4:0] ? 32'hbd6e2940 : _GEN_1968; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1970 = 5'h17 == _T_220[4:0] ? 32'hbf7e44de : _GEN_1969; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1971 = 5'h18 == _T_220[4:0] ? 32'h3f800000 : _GEN_1970; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1972 = 5'h19 == _T_220[4:0] ? 32'hbe92d7dc : _GEN_1971; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_1978 = 5'h4 == _T_220[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1979 = 5'h5 == _T_220[4:0] ? 32'hbee5c900 : _GEN_1978; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1980 = 5'h6 == _T_220[4:0] ? 32'h80800000 : _GEN_1979; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1981 = 5'h7 == _T_220[4:0] ? 32'hbee5c900 : _GEN_1980; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1982 = 5'h8 == _T_220[4:0] ? 32'hbf4d57f2 : _GEN_1981; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1983 = 5'h9 == _T_220[4:0] ? 32'h80800000 : _GEN_1982; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1984 = 5'ha == _T_220[4:0] ? 32'hbf248dba : _GEN_1983; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1985 = 5'hb == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1984; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1986 = 5'hc == _T_220[4:0] ? 32'h80800000 : _GEN_1985; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1987 = 5'hd == _T_220[4:0] ? 32'hbf4d57f2 : _GEN_1986; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1988 = 5'he == _T_220[4:0] ? 32'hbf753ecc : _GEN_1987; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1989 = 5'hf == _T_220[4:0] ? 32'h80800000 : _GEN_1988; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1990 = 5'h10 == _T_220[4:0] ? 32'hbf6b1034 : _GEN_1989; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1991 = 5'h11 == _T_220[4:0] ? 32'hbf3a3528 : _GEN_1990; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1992 = 5'h12 == _T_220[4:0] ? 32'h80800000 : _GEN_1991; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1993 = 5'h13 == _T_220[4:0] ? 32'hbf7c1c5c : _GEN_1992; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1994 = 5'h14 == _T_220[4:0] ? 32'hbeaf1d40 : _GEN_1993; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1995 = 5'h15 == _T_220[4:0] ? 32'h80800000 : _GEN_1994; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1996 = 5'h16 == _T_220[4:0] ? 32'hbf7f911e : _GEN_1995; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1997 = 5'h17 == _T_220[4:0] ? 32'h3dedc210 : _GEN_1996; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1998 = 5'h18 == _T_220[4:0] ? 32'h80800000 : _GEN_1997; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_1999 = 5'h19 == _T_220[4:0] ? 32'hbf753ecc : _GEN_1998; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2002 = 5'h1 == _T_220[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2003 = 5'h2 == _T_220[4:0] ? io_in_2_Im : _GEN_2002; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2004 = 5'h3 == _T_220[4:0] ? io_in_3_Im : _GEN_2003; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2005 = 5'h4 == _T_220[4:0] ? io_in_4_Im : _GEN_2004; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2006 = 5'h5 == _T_220[4:0] ? io_in_5_Im : _GEN_2005; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2007 = 5'h6 == _T_220[4:0] ? io_in_6_Im : _GEN_2006; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2008 = 5'h7 == _T_220[4:0] ? io_in_7_Im : _GEN_2007; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2009 = 5'h8 == _T_220[4:0] ? io_in_8_Im : _GEN_2008; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2010 = 5'h9 == _T_220[4:0] ? io_in_9_Im : _GEN_2009; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2011 = 5'ha == _T_220[4:0] ? io_in_10_Im : _GEN_2010; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2012 = 5'hb == _T_220[4:0] ? io_in_11_Im : _GEN_2011; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2013 = 5'hc == _T_220[4:0] ? io_in_12_Im : _GEN_2012; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2014 = 5'hd == _T_220[4:0] ? io_in_13_Im : _GEN_2013; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2015 = 5'he == _T_220[4:0] ? io_in_14_Im : _GEN_2014; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2016 = 5'hf == _T_220[4:0] ? io_in_15_Im : _GEN_2015; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2017 = 5'h10 == _T_220[4:0] ? io_in_16_Im : _GEN_2016; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2018 = 5'h11 == _T_220[4:0] ? io_in_17_Im : _GEN_2017; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2019 = 5'h12 == _T_220[4:0] ? io_in_18_Im : _GEN_2018; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2020 = 5'h13 == _T_220[4:0] ? io_in_19_Im : _GEN_2019; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2021 = 5'h14 == _T_220[4:0] ? io_in_20_Im : _GEN_2020; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2022 = 5'h15 == _T_220[4:0] ? io_in_21_Im : _GEN_2021; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2023 = 5'h16 == _T_220[4:0] ? io_in_22_Im : _GEN_2022; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2024 = 5'h17 == _T_220[4:0] ? io_in_23_Im : _GEN_2023; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2025 = 5'h18 == _T_220[4:0] ? io_in_24_Im : _GEN_2024; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2026 = 5'h19 == _T_220[4:0] ? io_in_25_Im : _GEN_2025; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2029 = 5'h1 == _T_220[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2030 = 5'h2 == _T_220[4:0] ? io_in_2_Re : _GEN_2029; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2031 = 5'h3 == _T_220[4:0] ? io_in_3_Re : _GEN_2030; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2032 = 5'h4 == _T_220[4:0] ? io_in_4_Re : _GEN_2031; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2033 = 5'h5 == _T_220[4:0] ? io_in_5_Re : _GEN_2032; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2034 = 5'h6 == _T_220[4:0] ? io_in_6_Re : _GEN_2033; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2035 = 5'h7 == _T_220[4:0] ? io_in_7_Re : _GEN_2034; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2036 = 5'h8 == _T_220[4:0] ? io_in_8_Re : _GEN_2035; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2037 = 5'h9 == _T_220[4:0] ? io_in_9_Re : _GEN_2036; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2038 = 5'ha == _T_220[4:0] ? io_in_10_Re : _GEN_2037; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2039 = 5'hb == _T_220[4:0] ? io_in_11_Re : _GEN_2038; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2040 = 5'hc == _T_220[4:0] ? io_in_12_Re : _GEN_2039; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2041 = 5'hd == _T_220[4:0] ? io_in_13_Re : _GEN_2040; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2042 = 5'he == _T_220[4:0] ? io_in_14_Re : _GEN_2041; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2043 = 5'hf == _T_220[4:0] ? io_in_15_Re : _GEN_2042; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2044 = 5'h10 == _T_220[4:0] ? io_in_16_Re : _GEN_2043; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2045 = 5'h11 == _T_220[4:0] ? io_in_17_Re : _GEN_2044; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2046 = 5'h12 == _T_220[4:0] ? io_in_18_Re : _GEN_2045; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2047 = 5'h13 == _T_220[4:0] ? io_in_19_Re : _GEN_2046; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2048 = 5'h14 == _T_220[4:0] ? io_in_20_Re : _GEN_2047; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2049 = 5'h15 == _T_220[4:0] ? io_in_21_Re : _GEN_2048; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2050 = 5'h16 == _T_220[4:0] ? io_in_22_Re : _GEN_2049; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2051 = 5'h17 == _T_220[4:0] ? io_in_23_Re : _GEN_2050; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2052 = 5'h18 == _T_220[4:0] ? io_in_24_Re : _GEN_2051; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2053 = 5'h19 == _T_220[4:0] ? io_in_25_Re : _GEN_2052; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_232 = _T_2 + 37'h13; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2059 = 5'h4 == _T_232[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2060 = 5'h5 == _T_232[4:0] ? 32'h3f64c51a : _GEN_2059; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2061 = 5'h6 == _T_232[4:0] ? 32'h3f800000 : _GEN_2060; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2062 = 5'h7 == _T_232[4:0] ? 32'h3f64c51a : _GEN_2061; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2063 = 5'h8 == _T_232[4:0] ? 32'h3f18df62 : _GEN_2062; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2064 = 5'h9 == _T_232[4:0] ? 32'h3f800000 : _GEN_2063; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2065 = 5'ha == _T_232[4:0] ? 32'h3f441b7c : _GEN_2064; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2066 = 5'hb == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2065; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2067 = 5'hc == _T_232[4:0] ? 32'h3f800000 : _GEN_2066; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2068 = 5'hd == _T_232[4:0] ? 32'h3f18df62 : _GEN_2067; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2069 = 5'he == _T_232[4:0] ? 32'hbe92d7dc : _GEN_2068; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2070 = 5'hf == _T_232[4:0] ? 32'h3f800000 : _GEN_2069; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2071 = 5'h10 == _T_232[4:0] ? 32'h3ecacaf4 : _GEN_2070; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2072 = 5'h11 == _T_232[4:0] ? 32'hbf2fad88 : _GEN_2071; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2073 = 5'h12 == _T_232[4:0] ? 32'h3f800000 : _GEN_2072; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2074 = 5'h13 == _T_232[4:0] ? 32'h3e31d0d0 : _GEN_2073; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2075 = 5'h14 == _T_232[4:0] ? 32'hbf708fb2 : _GEN_2074; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2076 = 5'h15 == _T_232[4:0] ? 32'h3f800000 : _GEN_2075; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2077 = 5'h16 == _T_232[4:0] ? 32'hbd6e2940 : _GEN_2076; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2078 = 5'h17 == _T_232[4:0] ? 32'hbf7e44de : _GEN_2077; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2079 = 5'h18 == _T_232[4:0] ? 32'h3f800000 : _GEN_2078; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2080 = 5'h19 == _T_232[4:0] ? 32'hbe92d7dc : _GEN_2079; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2086 = 5'h4 == _T_232[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2087 = 5'h5 == _T_232[4:0] ? 32'hbee5c900 : _GEN_2086; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2088 = 5'h6 == _T_232[4:0] ? 32'h80800000 : _GEN_2087; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2089 = 5'h7 == _T_232[4:0] ? 32'hbee5c900 : _GEN_2088; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2090 = 5'h8 == _T_232[4:0] ? 32'hbf4d57f2 : _GEN_2089; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2091 = 5'h9 == _T_232[4:0] ? 32'h80800000 : _GEN_2090; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2092 = 5'ha == _T_232[4:0] ? 32'hbf248dba : _GEN_2091; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2093 = 5'hb == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2092; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2094 = 5'hc == _T_232[4:0] ? 32'h80800000 : _GEN_2093; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2095 = 5'hd == _T_232[4:0] ? 32'hbf4d57f2 : _GEN_2094; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2096 = 5'he == _T_232[4:0] ? 32'hbf753ecc : _GEN_2095; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2097 = 5'hf == _T_232[4:0] ? 32'h80800000 : _GEN_2096; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2098 = 5'h10 == _T_232[4:0] ? 32'hbf6b1034 : _GEN_2097; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2099 = 5'h11 == _T_232[4:0] ? 32'hbf3a3528 : _GEN_2098; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2100 = 5'h12 == _T_232[4:0] ? 32'h80800000 : _GEN_2099; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2101 = 5'h13 == _T_232[4:0] ? 32'hbf7c1c5c : _GEN_2100; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2102 = 5'h14 == _T_232[4:0] ? 32'hbeaf1d40 : _GEN_2101; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2103 = 5'h15 == _T_232[4:0] ? 32'h80800000 : _GEN_2102; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2104 = 5'h16 == _T_232[4:0] ? 32'hbf7f911e : _GEN_2103; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2105 = 5'h17 == _T_232[4:0] ? 32'h3dedc210 : _GEN_2104; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2106 = 5'h18 == _T_232[4:0] ? 32'h80800000 : _GEN_2105; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2107 = 5'h19 == _T_232[4:0] ? 32'hbf753ecc : _GEN_2106; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2110 = 5'h1 == _T_232[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2111 = 5'h2 == _T_232[4:0] ? io_in_2_Im : _GEN_2110; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2112 = 5'h3 == _T_232[4:0] ? io_in_3_Im : _GEN_2111; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2113 = 5'h4 == _T_232[4:0] ? io_in_4_Im : _GEN_2112; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2114 = 5'h5 == _T_232[4:0] ? io_in_5_Im : _GEN_2113; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2115 = 5'h6 == _T_232[4:0] ? io_in_6_Im : _GEN_2114; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2116 = 5'h7 == _T_232[4:0] ? io_in_7_Im : _GEN_2115; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2117 = 5'h8 == _T_232[4:0] ? io_in_8_Im : _GEN_2116; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2118 = 5'h9 == _T_232[4:0] ? io_in_9_Im : _GEN_2117; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2119 = 5'ha == _T_232[4:0] ? io_in_10_Im : _GEN_2118; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2120 = 5'hb == _T_232[4:0] ? io_in_11_Im : _GEN_2119; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2121 = 5'hc == _T_232[4:0] ? io_in_12_Im : _GEN_2120; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2122 = 5'hd == _T_232[4:0] ? io_in_13_Im : _GEN_2121; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2123 = 5'he == _T_232[4:0] ? io_in_14_Im : _GEN_2122; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2124 = 5'hf == _T_232[4:0] ? io_in_15_Im : _GEN_2123; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2125 = 5'h10 == _T_232[4:0] ? io_in_16_Im : _GEN_2124; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2126 = 5'h11 == _T_232[4:0] ? io_in_17_Im : _GEN_2125; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2127 = 5'h12 == _T_232[4:0] ? io_in_18_Im : _GEN_2126; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2128 = 5'h13 == _T_232[4:0] ? io_in_19_Im : _GEN_2127; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2129 = 5'h14 == _T_232[4:0] ? io_in_20_Im : _GEN_2128; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2130 = 5'h15 == _T_232[4:0] ? io_in_21_Im : _GEN_2129; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2131 = 5'h16 == _T_232[4:0] ? io_in_22_Im : _GEN_2130; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2132 = 5'h17 == _T_232[4:0] ? io_in_23_Im : _GEN_2131; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2133 = 5'h18 == _T_232[4:0] ? io_in_24_Im : _GEN_2132; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2134 = 5'h19 == _T_232[4:0] ? io_in_25_Im : _GEN_2133; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2137 = 5'h1 == _T_232[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2138 = 5'h2 == _T_232[4:0] ? io_in_2_Re : _GEN_2137; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2139 = 5'h3 == _T_232[4:0] ? io_in_3_Re : _GEN_2138; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2140 = 5'h4 == _T_232[4:0] ? io_in_4_Re : _GEN_2139; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2141 = 5'h5 == _T_232[4:0] ? io_in_5_Re : _GEN_2140; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2142 = 5'h6 == _T_232[4:0] ? io_in_6_Re : _GEN_2141; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2143 = 5'h7 == _T_232[4:0] ? io_in_7_Re : _GEN_2142; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2144 = 5'h8 == _T_232[4:0] ? io_in_8_Re : _GEN_2143; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2145 = 5'h9 == _T_232[4:0] ? io_in_9_Re : _GEN_2144; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2146 = 5'ha == _T_232[4:0] ? io_in_10_Re : _GEN_2145; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2147 = 5'hb == _T_232[4:0] ? io_in_11_Re : _GEN_2146; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2148 = 5'hc == _T_232[4:0] ? io_in_12_Re : _GEN_2147; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2149 = 5'hd == _T_232[4:0] ? io_in_13_Re : _GEN_2148; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2150 = 5'he == _T_232[4:0] ? io_in_14_Re : _GEN_2149; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2151 = 5'hf == _T_232[4:0] ? io_in_15_Re : _GEN_2150; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2152 = 5'h10 == _T_232[4:0] ? io_in_16_Re : _GEN_2151; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2153 = 5'h11 == _T_232[4:0] ? io_in_17_Re : _GEN_2152; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2154 = 5'h12 == _T_232[4:0] ? io_in_18_Re : _GEN_2153; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2155 = 5'h13 == _T_232[4:0] ? io_in_19_Re : _GEN_2154; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2156 = 5'h14 == _T_232[4:0] ? io_in_20_Re : _GEN_2155; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2157 = 5'h15 == _T_232[4:0] ? io_in_21_Re : _GEN_2156; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2158 = 5'h16 == _T_232[4:0] ? io_in_22_Re : _GEN_2157; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2159 = 5'h17 == _T_232[4:0] ? io_in_23_Re : _GEN_2158; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2160 = 5'h18 == _T_232[4:0] ? io_in_24_Re : _GEN_2159; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2161 = 5'h19 == _T_232[4:0] ? io_in_25_Re : _GEN_2160; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_244 = _T_2 + 37'h14; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2167 = 5'h4 == _T_244[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2168 = 5'h5 == _T_244[4:0] ? 32'h3f64c51a : _GEN_2167; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2169 = 5'h6 == _T_244[4:0] ? 32'h3f800000 : _GEN_2168; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2170 = 5'h7 == _T_244[4:0] ? 32'h3f64c51a : _GEN_2169; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2171 = 5'h8 == _T_244[4:0] ? 32'h3f18df62 : _GEN_2170; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2172 = 5'h9 == _T_244[4:0] ? 32'h3f800000 : _GEN_2171; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2173 = 5'ha == _T_244[4:0] ? 32'h3f441b7c : _GEN_2172; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2174 = 5'hb == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2173; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2175 = 5'hc == _T_244[4:0] ? 32'h3f800000 : _GEN_2174; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2176 = 5'hd == _T_244[4:0] ? 32'h3f18df62 : _GEN_2175; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2177 = 5'he == _T_244[4:0] ? 32'hbe92d7dc : _GEN_2176; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2178 = 5'hf == _T_244[4:0] ? 32'h3f800000 : _GEN_2177; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2179 = 5'h10 == _T_244[4:0] ? 32'h3ecacaf4 : _GEN_2178; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2180 = 5'h11 == _T_244[4:0] ? 32'hbf2fad88 : _GEN_2179; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2181 = 5'h12 == _T_244[4:0] ? 32'h3f800000 : _GEN_2180; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2182 = 5'h13 == _T_244[4:0] ? 32'h3e31d0d0 : _GEN_2181; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2183 = 5'h14 == _T_244[4:0] ? 32'hbf708fb2 : _GEN_2182; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2184 = 5'h15 == _T_244[4:0] ? 32'h3f800000 : _GEN_2183; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2185 = 5'h16 == _T_244[4:0] ? 32'hbd6e2940 : _GEN_2184; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2186 = 5'h17 == _T_244[4:0] ? 32'hbf7e44de : _GEN_2185; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2187 = 5'h18 == _T_244[4:0] ? 32'h3f800000 : _GEN_2186; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2188 = 5'h19 == _T_244[4:0] ? 32'hbe92d7dc : _GEN_2187; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2194 = 5'h4 == _T_244[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2195 = 5'h5 == _T_244[4:0] ? 32'hbee5c900 : _GEN_2194; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2196 = 5'h6 == _T_244[4:0] ? 32'h80800000 : _GEN_2195; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2197 = 5'h7 == _T_244[4:0] ? 32'hbee5c900 : _GEN_2196; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2198 = 5'h8 == _T_244[4:0] ? 32'hbf4d57f2 : _GEN_2197; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2199 = 5'h9 == _T_244[4:0] ? 32'h80800000 : _GEN_2198; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2200 = 5'ha == _T_244[4:0] ? 32'hbf248dba : _GEN_2199; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2201 = 5'hb == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2200; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2202 = 5'hc == _T_244[4:0] ? 32'h80800000 : _GEN_2201; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2203 = 5'hd == _T_244[4:0] ? 32'hbf4d57f2 : _GEN_2202; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2204 = 5'he == _T_244[4:0] ? 32'hbf753ecc : _GEN_2203; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2205 = 5'hf == _T_244[4:0] ? 32'h80800000 : _GEN_2204; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2206 = 5'h10 == _T_244[4:0] ? 32'hbf6b1034 : _GEN_2205; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2207 = 5'h11 == _T_244[4:0] ? 32'hbf3a3528 : _GEN_2206; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2208 = 5'h12 == _T_244[4:0] ? 32'h80800000 : _GEN_2207; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2209 = 5'h13 == _T_244[4:0] ? 32'hbf7c1c5c : _GEN_2208; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2210 = 5'h14 == _T_244[4:0] ? 32'hbeaf1d40 : _GEN_2209; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2211 = 5'h15 == _T_244[4:0] ? 32'h80800000 : _GEN_2210; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2212 = 5'h16 == _T_244[4:0] ? 32'hbf7f911e : _GEN_2211; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2213 = 5'h17 == _T_244[4:0] ? 32'h3dedc210 : _GEN_2212; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2214 = 5'h18 == _T_244[4:0] ? 32'h80800000 : _GEN_2213; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2215 = 5'h19 == _T_244[4:0] ? 32'hbf753ecc : _GEN_2214; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2218 = 5'h1 == _T_244[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2219 = 5'h2 == _T_244[4:0] ? io_in_2_Im : _GEN_2218; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2220 = 5'h3 == _T_244[4:0] ? io_in_3_Im : _GEN_2219; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2221 = 5'h4 == _T_244[4:0] ? io_in_4_Im : _GEN_2220; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2222 = 5'h5 == _T_244[4:0] ? io_in_5_Im : _GEN_2221; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2223 = 5'h6 == _T_244[4:0] ? io_in_6_Im : _GEN_2222; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2224 = 5'h7 == _T_244[4:0] ? io_in_7_Im : _GEN_2223; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2225 = 5'h8 == _T_244[4:0] ? io_in_8_Im : _GEN_2224; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2226 = 5'h9 == _T_244[4:0] ? io_in_9_Im : _GEN_2225; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2227 = 5'ha == _T_244[4:0] ? io_in_10_Im : _GEN_2226; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2228 = 5'hb == _T_244[4:0] ? io_in_11_Im : _GEN_2227; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2229 = 5'hc == _T_244[4:0] ? io_in_12_Im : _GEN_2228; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2230 = 5'hd == _T_244[4:0] ? io_in_13_Im : _GEN_2229; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2231 = 5'he == _T_244[4:0] ? io_in_14_Im : _GEN_2230; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2232 = 5'hf == _T_244[4:0] ? io_in_15_Im : _GEN_2231; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2233 = 5'h10 == _T_244[4:0] ? io_in_16_Im : _GEN_2232; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2234 = 5'h11 == _T_244[4:0] ? io_in_17_Im : _GEN_2233; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2235 = 5'h12 == _T_244[4:0] ? io_in_18_Im : _GEN_2234; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2236 = 5'h13 == _T_244[4:0] ? io_in_19_Im : _GEN_2235; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2237 = 5'h14 == _T_244[4:0] ? io_in_20_Im : _GEN_2236; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2238 = 5'h15 == _T_244[4:0] ? io_in_21_Im : _GEN_2237; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2239 = 5'h16 == _T_244[4:0] ? io_in_22_Im : _GEN_2238; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2240 = 5'h17 == _T_244[4:0] ? io_in_23_Im : _GEN_2239; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2241 = 5'h18 == _T_244[4:0] ? io_in_24_Im : _GEN_2240; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2242 = 5'h19 == _T_244[4:0] ? io_in_25_Im : _GEN_2241; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2245 = 5'h1 == _T_244[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2246 = 5'h2 == _T_244[4:0] ? io_in_2_Re : _GEN_2245; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2247 = 5'h3 == _T_244[4:0] ? io_in_3_Re : _GEN_2246; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2248 = 5'h4 == _T_244[4:0] ? io_in_4_Re : _GEN_2247; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2249 = 5'h5 == _T_244[4:0] ? io_in_5_Re : _GEN_2248; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2250 = 5'h6 == _T_244[4:0] ? io_in_6_Re : _GEN_2249; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2251 = 5'h7 == _T_244[4:0] ? io_in_7_Re : _GEN_2250; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2252 = 5'h8 == _T_244[4:0] ? io_in_8_Re : _GEN_2251; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2253 = 5'h9 == _T_244[4:0] ? io_in_9_Re : _GEN_2252; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2254 = 5'ha == _T_244[4:0] ? io_in_10_Re : _GEN_2253; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2255 = 5'hb == _T_244[4:0] ? io_in_11_Re : _GEN_2254; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2256 = 5'hc == _T_244[4:0] ? io_in_12_Re : _GEN_2255; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2257 = 5'hd == _T_244[4:0] ? io_in_13_Re : _GEN_2256; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2258 = 5'he == _T_244[4:0] ? io_in_14_Re : _GEN_2257; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2259 = 5'hf == _T_244[4:0] ? io_in_15_Re : _GEN_2258; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2260 = 5'h10 == _T_244[4:0] ? io_in_16_Re : _GEN_2259; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2261 = 5'h11 == _T_244[4:0] ? io_in_17_Re : _GEN_2260; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2262 = 5'h12 == _T_244[4:0] ? io_in_18_Re : _GEN_2261; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2263 = 5'h13 == _T_244[4:0] ? io_in_19_Re : _GEN_2262; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2264 = 5'h14 == _T_244[4:0] ? io_in_20_Re : _GEN_2263; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2265 = 5'h15 == _T_244[4:0] ? io_in_21_Re : _GEN_2264; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2266 = 5'h16 == _T_244[4:0] ? io_in_22_Re : _GEN_2265; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2267 = 5'h17 == _T_244[4:0] ? io_in_23_Re : _GEN_2266; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2268 = 5'h18 == _T_244[4:0] ? io_in_24_Re : _GEN_2267; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2269 = 5'h19 == _T_244[4:0] ? io_in_25_Re : _GEN_2268; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_256 = _T_2 + 37'h15; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2275 = 5'h4 == _T_256[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2276 = 5'h5 == _T_256[4:0] ? 32'h3f64c51a : _GEN_2275; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2277 = 5'h6 == _T_256[4:0] ? 32'h3f800000 : _GEN_2276; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2278 = 5'h7 == _T_256[4:0] ? 32'h3f64c51a : _GEN_2277; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2279 = 5'h8 == _T_256[4:0] ? 32'h3f18df62 : _GEN_2278; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2280 = 5'h9 == _T_256[4:0] ? 32'h3f800000 : _GEN_2279; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2281 = 5'ha == _T_256[4:0] ? 32'h3f441b7c : _GEN_2280; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2282 = 5'hb == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2281; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2283 = 5'hc == _T_256[4:0] ? 32'h3f800000 : _GEN_2282; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2284 = 5'hd == _T_256[4:0] ? 32'h3f18df62 : _GEN_2283; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2285 = 5'he == _T_256[4:0] ? 32'hbe92d7dc : _GEN_2284; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2286 = 5'hf == _T_256[4:0] ? 32'h3f800000 : _GEN_2285; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2287 = 5'h10 == _T_256[4:0] ? 32'h3ecacaf4 : _GEN_2286; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2288 = 5'h11 == _T_256[4:0] ? 32'hbf2fad88 : _GEN_2287; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2289 = 5'h12 == _T_256[4:0] ? 32'h3f800000 : _GEN_2288; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2290 = 5'h13 == _T_256[4:0] ? 32'h3e31d0d0 : _GEN_2289; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2291 = 5'h14 == _T_256[4:0] ? 32'hbf708fb2 : _GEN_2290; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2292 = 5'h15 == _T_256[4:0] ? 32'h3f800000 : _GEN_2291; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2293 = 5'h16 == _T_256[4:0] ? 32'hbd6e2940 : _GEN_2292; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2294 = 5'h17 == _T_256[4:0] ? 32'hbf7e44de : _GEN_2293; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2295 = 5'h18 == _T_256[4:0] ? 32'h3f800000 : _GEN_2294; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2296 = 5'h19 == _T_256[4:0] ? 32'hbe92d7dc : _GEN_2295; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2302 = 5'h4 == _T_256[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2303 = 5'h5 == _T_256[4:0] ? 32'hbee5c900 : _GEN_2302; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2304 = 5'h6 == _T_256[4:0] ? 32'h80800000 : _GEN_2303; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2305 = 5'h7 == _T_256[4:0] ? 32'hbee5c900 : _GEN_2304; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2306 = 5'h8 == _T_256[4:0] ? 32'hbf4d57f2 : _GEN_2305; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2307 = 5'h9 == _T_256[4:0] ? 32'h80800000 : _GEN_2306; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2308 = 5'ha == _T_256[4:0] ? 32'hbf248dba : _GEN_2307; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2309 = 5'hb == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2308; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2310 = 5'hc == _T_256[4:0] ? 32'h80800000 : _GEN_2309; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2311 = 5'hd == _T_256[4:0] ? 32'hbf4d57f2 : _GEN_2310; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2312 = 5'he == _T_256[4:0] ? 32'hbf753ecc : _GEN_2311; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2313 = 5'hf == _T_256[4:0] ? 32'h80800000 : _GEN_2312; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2314 = 5'h10 == _T_256[4:0] ? 32'hbf6b1034 : _GEN_2313; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2315 = 5'h11 == _T_256[4:0] ? 32'hbf3a3528 : _GEN_2314; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2316 = 5'h12 == _T_256[4:0] ? 32'h80800000 : _GEN_2315; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2317 = 5'h13 == _T_256[4:0] ? 32'hbf7c1c5c : _GEN_2316; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2318 = 5'h14 == _T_256[4:0] ? 32'hbeaf1d40 : _GEN_2317; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2319 = 5'h15 == _T_256[4:0] ? 32'h80800000 : _GEN_2318; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2320 = 5'h16 == _T_256[4:0] ? 32'hbf7f911e : _GEN_2319; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2321 = 5'h17 == _T_256[4:0] ? 32'h3dedc210 : _GEN_2320; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2322 = 5'h18 == _T_256[4:0] ? 32'h80800000 : _GEN_2321; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2323 = 5'h19 == _T_256[4:0] ? 32'hbf753ecc : _GEN_2322; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2326 = 5'h1 == _T_256[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2327 = 5'h2 == _T_256[4:0] ? io_in_2_Im : _GEN_2326; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2328 = 5'h3 == _T_256[4:0] ? io_in_3_Im : _GEN_2327; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2329 = 5'h4 == _T_256[4:0] ? io_in_4_Im : _GEN_2328; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2330 = 5'h5 == _T_256[4:0] ? io_in_5_Im : _GEN_2329; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2331 = 5'h6 == _T_256[4:0] ? io_in_6_Im : _GEN_2330; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2332 = 5'h7 == _T_256[4:0] ? io_in_7_Im : _GEN_2331; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2333 = 5'h8 == _T_256[4:0] ? io_in_8_Im : _GEN_2332; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2334 = 5'h9 == _T_256[4:0] ? io_in_9_Im : _GEN_2333; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2335 = 5'ha == _T_256[4:0] ? io_in_10_Im : _GEN_2334; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2336 = 5'hb == _T_256[4:0] ? io_in_11_Im : _GEN_2335; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2337 = 5'hc == _T_256[4:0] ? io_in_12_Im : _GEN_2336; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2338 = 5'hd == _T_256[4:0] ? io_in_13_Im : _GEN_2337; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2339 = 5'he == _T_256[4:0] ? io_in_14_Im : _GEN_2338; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2340 = 5'hf == _T_256[4:0] ? io_in_15_Im : _GEN_2339; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2341 = 5'h10 == _T_256[4:0] ? io_in_16_Im : _GEN_2340; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2342 = 5'h11 == _T_256[4:0] ? io_in_17_Im : _GEN_2341; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2343 = 5'h12 == _T_256[4:0] ? io_in_18_Im : _GEN_2342; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2344 = 5'h13 == _T_256[4:0] ? io_in_19_Im : _GEN_2343; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2345 = 5'h14 == _T_256[4:0] ? io_in_20_Im : _GEN_2344; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2346 = 5'h15 == _T_256[4:0] ? io_in_21_Im : _GEN_2345; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2347 = 5'h16 == _T_256[4:0] ? io_in_22_Im : _GEN_2346; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2348 = 5'h17 == _T_256[4:0] ? io_in_23_Im : _GEN_2347; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2349 = 5'h18 == _T_256[4:0] ? io_in_24_Im : _GEN_2348; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2350 = 5'h19 == _T_256[4:0] ? io_in_25_Im : _GEN_2349; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2353 = 5'h1 == _T_256[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2354 = 5'h2 == _T_256[4:0] ? io_in_2_Re : _GEN_2353; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2355 = 5'h3 == _T_256[4:0] ? io_in_3_Re : _GEN_2354; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2356 = 5'h4 == _T_256[4:0] ? io_in_4_Re : _GEN_2355; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2357 = 5'h5 == _T_256[4:0] ? io_in_5_Re : _GEN_2356; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2358 = 5'h6 == _T_256[4:0] ? io_in_6_Re : _GEN_2357; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2359 = 5'h7 == _T_256[4:0] ? io_in_7_Re : _GEN_2358; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2360 = 5'h8 == _T_256[4:0] ? io_in_8_Re : _GEN_2359; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2361 = 5'h9 == _T_256[4:0] ? io_in_9_Re : _GEN_2360; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2362 = 5'ha == _T_256[4:0] ? io_in_10_Re : _GEN_2361; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2363 = 5'hb == _T_256[4:0] ? io_in_11_Re : _GEN_2362; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2364 = 5'hc == _T_256[4:0] ? io_in_12_Re : _GEN_2363; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2365 = 5'hd == _T_256[4:0] ? io_in_13_Re : _GEN_2364; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2366 = 5'he == _T_256[4:0] ? io_in_14_Re : _GEN_2365; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2367 = 5'hf == _T_256[4:0] ? io_in_15_Re : _GEN_2366; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2368 = 5'h10 == _T_256[4:0] ? io_in_16_Re : _GEN_2367; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2369 = 5'h11 == _T_256[4:0] ? io_in_17_Re : _GEN_2368; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2370 = 5'h12 == _T_256[4:0] ? io_in_18_Re : _GEN_2369; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2371 = 5'h13 == _T_256[4:0] ? io_in_19_Re : _GEN_2370; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2372 = 5'h14 == _T_256[4:0] ? io_in_20_Re : _GEN_2371; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2373 = 5'h15 == _T_256[4:0] ? io_in_21_Re : _GEN_2372; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2374 = 5'h16 == _T_256[4:0] ? io_in_22_Re : _GEN_2373; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2375 = 5'h17 == _T_256[4:0] ? io_in_23_Re : _GEN_2374; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2376 = 5'h18 == _T_256[4:0] ? io_in_24_Re : _GEN_2375; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2377 = 5'h19 == _T_256[4:0] ? io_in_25_Re : _GEN_2376; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_268 = _T_2 + 37'h16; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2383 = 5'h4 == _T_268[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2384 = 5'h5 == _T_268[4:0] ? 32'h3f64c51a : _GEN_2383; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2385 = 5'h6 == _T_268[4:0] ? 32'h3f800000 : _GEN_2384; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2386 = 5'h7 == _T_268[4:0] ? 32'h3f64c51a : _GEN_2385; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2387 = 5'h8 == _T_268[4:0] ? 32'h3f18df62 : _GEN_2386; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2388 = 5'h9 == _T_268[4:0] ? 32'h3f800000 : _GEN_2387; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2389 = 5'ha == _T_268[4:0] ? 32'h3f441b7c : _GEN_2388; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2390 = 5'hb == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2389; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2391 = 5'hc == _T_268[4:0] ? 32'h3f800000 : _GEN_2390; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2392 = 5'hd == _T_268[4:0] ? 32'h3f18df62 : _GEN_2391; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2393 = 5'he == _T_268[4:0] ? 32'hbe92d7dc : _GEN_2392; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2394 = 5'hf == _T_268[4:0] ? 32'h3f800000 : _GEN_2393; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2395 = 5'h10 == _T_268[4:0] ? 32'h3ecacaf4 : _GEN_2394; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2396 = 5'h11 == _T_268[4:0] ? 32'hbf2fad88 : _GEN_2395; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2397 = 5'h12 == _T_268[4:0] ? 32'h3f800000 : _GEN_2396; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2398 = 5'h13 == _T_268[4:0] ? 32'h3e31d0d0 : _GEN_2397; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2399 = 5'h14 == _T_268[4:0] ? 32'hbf708fb2 : _GEN_2398; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2400 = 5'h15 == _T_268[4:0] ? 32'h3f800000 : _GEN_2399; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2401 = 5'h16 == _T_268[4:0] ? 32'hbd6e2940 : _GEN_2400; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2402 = 5'h17 == _T_268[4:0] ? 32'hbf7e44de : _GEN_2401; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2403 = 5'h18 == _T_268[4:0] ? 32'h3f800000 : _GEN_2402; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2404 = 5'h19 == _T_268[4:0] ? 32'hbe92d7dc : _GEN_2403; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2410 = 5'h4 == _T_268[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2411 = 5'h5 == _T_268[4:0] ? 32'hbee5c900 : _GEN_2410; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2412 = 5'h6 == _T_268[4:0] ? 32'h80800000 : _GEN_2411; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2413 = 5'h7 == _T_268[4:0] ? 32'hbee5c900 : _GEN_2412; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2414 = 5'h8 == _T_268[4:0] ? 32'hbf4d57f2 : _GEN_2413; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2415 = 5'h9 == _T_268[4:0] ? 32'h80800000 : _GEN_2414; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2416 = 5'ha == _T_268[4:0] ? 32'hbf248dba : _GEN_2415; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2417 = 5'hb == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2416; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2418 = 5'hc == _T_268[4:0] ? 32'h80800000 : _GEN_2417; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2419 = 5'hd == _T_268[4:0] ? 32'hbf4d57f2 : _GEN_2418; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2420 = 5'he == _T_268[4:0] ? 32'hbf753ecc : _GEN_2419; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2421 = 5'hf == _T_268[4:0] ? 32'h80800000 : _GEN_2420; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2422 = 5'h10 == _T_268[4:0] ? 32'hbf6b1034 : _GEN_2421; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2423 = 5'h11 == _T_268[4:0] ? 32'hbf3a3528 : _GEN_2422; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2424 = 5'h12 == _T_268[4:0] ? 32'h80800000 : _GEN_2423; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2425 = 5'h13 == _T_268[4:0] ? 32'hbf7c1c5c : _GEN_2424; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2426 = 5'h14 == _T_268[4:0] ? 32'hbeaf1d40 : _GEN_2425; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2427 = 5'h15 == _T_268[4:0] ? 32'h80800000 : _GEN_2426; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2428 = 5'h16 == _T_268[4:0] ? 32'hbf7f911e : _GEN_2427; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2429 = 5'h17 == _T_268[4:0] ? 32'h3dedc210 : _GEN_2428; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2430 = 5'h18 == _T_268[4:0] ? 32'h80800000 : _GEN_2429; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2431 = 5'h19 == _T_268[4:0] ? 32'hbf753ecc : _GEN_2430; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2434 = 5'h1 == _T_268[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2435 = 5'h2 == _T_268[4:0] ? io_in_2_Im : _GEN_2434; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2436 = 5'h3 == _T_268[4:0] ? io_in_3_Im : _GEN_2435; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2437 = 5'h4 == _T_268[4:0] ? io_in_4_Im : _GEN_2436; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2438 = 5'h5 == _T_268[4:0] ? io_in_5_Im : _GEN_2437; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2439 = 5'h6 == _T_268[4:0] ? io_in_6_Im : _GEN_2438; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2440 = 5'h7 == _T_268[4:0] ? io_in_7_Im : _GEN_2439; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2441 = 5'h8 == _T_268[4:0] ? io_in_8_Im : _GEN_2440; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2442 = 5'h9 == _T_268[4:0] ? io_in_9_Im : _GEN_2441; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2443 = 5'ha == _T_268[4:0] ? io_in_10_Im : _GEN_2442; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2444 = 5'hb == _T_268[4:0] ? io_in_11_Im : _GEN_2443; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2445 = 5'hc == _T_268[4:0] ? io_in_12_Im : _GEN_2444; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2446 = 5'hd == _T_268[4:0] ? io_in_13_Im : _GEN_2445; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2447 = 5'he == _T_268[4:0] ? io_in_14_Im : _GEN_2446; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2448 = 5'hf == _T_268[4:0] ? io_in_15_Im : _GEN_2447; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2449 = 5'h10 == _T_268[4:0] ? io_in_16_Im : _GEN_2448; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2450 = 5'h11 == _T_268[4:0] ? io_in_17_Im : _GEN_2449; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2451 = 5'h12 == _T_268[4:0] ? io_in_18_Im : _GEN_2450; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2452 = 5'h13 == _T_268[4:0] ? io_in_19_Im : _GEN_2451; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2453 = 5'h14 == _T_268[4:0] ? io_in_20_Im : _GEN_2452; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2454 = 5'h15 == _T_268[4:0] ? io_in_21_Im : _GEN_2453; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2455 = 5'h16 == _T_268[4:0] ? io_in_22_Im : _GEN_2454; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2456 = 5'h17 == _T_268[4:0] ? io_in_23_Im : _GEN_2455; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2457 = 5'h18 == _T_268[4:0] ? io_in_24_Im : _GEN_2456; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2458 = 5'h19 == _T_268[4:0] ? io_in_25_Im : _GEN_2457; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2461 = 5'h1 == _T_268[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2462 = 5'h2 == _T_268[4:0] ? io_in_2_Re : _GEN_2461; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2463 = 5'h3 == _T_268[4:0] ? io_in_3_Re : _GEN_2462; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2464 = 5'h4 == _T_268[4:0] ? io_in_4_Re : _GEN_2463; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2465 = 5'h5 == _T_268[4:0] ? io_in_5_Re : _GEN_2464; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2466 = 5'h6 == _T_268[4:0] ? io_in_6_Re : _GEN_2465; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2467 = 5'h7 == _T_268[4:0] ? io_in_7_Re : _GEN_2466; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2468 = 5'h8 == _T_268[4:0] ? io_in_8_Re : _GEN_2467; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2469 = 5'h9 == _T_268[4:0] ? io_in_9_Re : _GEN_2468; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2470 = 5'ha == _T_268[4:0] ? io_in_10_Re : _GEN_2469; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2471 = 5'hb == _T_268[4:0] ? io_in_11_Re : _GEN_2470; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2472 = 5'hc == _T_268[4:0] ? io_in_12_Re : _GEN_2471; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2473 = 5'hd == _T_268[4:0] ? io_in_13_Re : _GEN_2472; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2474 = 5'he == _T_268[4:0] ? io_in_14_Re : _GEN_2473; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2475 = 5'hf == _T_268[4:0] ? io_in_15_Re : _GEN_2474; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2476 = 5'h10 == _T_268[4:0] ? io_in_16_Re : _GEN_2475; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2477 = 5'h11 == _T_268[4:0] ? io_in_17_Re : _GEN_2476; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2478 = 5'h12 == _T_268[4:0] ? io_in_18_Re : _GEN_2477; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2479 = 5'h13 == _T_268[4:0] ? io_in_19_Re : _GEN_2478; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2480 = 5'h14 == _T_268[4:0] ? io_in_20_Re : _GEN_2479; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2481 = 5'h15 == _T_268[4:0] ? io_in_21_Re : _GEN_2480; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2482 = 5'h16 == _T_268[4:0] ? io_in_22_Re : _GEN_2481; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2483 = 5'h17 == _T_268[4:0] ? io_in_23_Re : _GEN_2482; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2484 = 5'h18 == _T_268[4:0] ? io_in_24_Re : _GEN_2483; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2485 = 5'h19 == _T_268[4:0] ? io_in_25_Re : _GEN_2484; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_280 = _T_2 + 37'h17; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2491 = 5'h4 == _T_280[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2492 = 5'h5 == _T_280[4:0] ? 32'h3f64c51a : _GEN_2491; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2493 = 5'h6 == _T_280[4:0] ? 32'h3f800000 : _GEN_2492; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2494 = 5'h7 == _T_280[4:0] ? 32'h3f64c51a : _GEN_2493; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2495 = 5'h8 == _T_280[4:0] ? 32'h3f18df62 : _GEN_2494; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2496 = 5'h9 == _T_280[4:0] ? 32'h3f800000 : _GEN_2495; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2497 = 5'ha == _T_280[4:0] ? 32'h3f441b7c : _GEN_2496; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2498 = 5'hb == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2497; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2499 = 5'hc == _T_280[4:0] ? 32'h3f800000 : _GEN_2498; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2500 = 5'hd == _T_280[4:0] ? 32'h3f18df62 : _GEN_2499; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2501 = 5'he == _T_280[4:0] ? 32'hbe92d7dc : _GEN_2500; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2502 = 5'hf == _T_280[4:0] ? 32'h3f800000 : _GEN_2501; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2503 = 5'h10 == _T_280[4:0] ? 32'h3ecacaf4 : _GEN_2502; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2504 = 5'h11 == _T_280[4:0] ? 32'hbf2fad88 : _GEN_2503; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2505 = 5'h12 == _T_280[4:0] ? 32'h3f800000 : _GEN_2504; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2506 = 5'h13 == _T_280[4:0] ? 32'h3e31d0d0 : _GEN_2505; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2507 = 5'h14 == _T_280[4:0] ? 32'hbf708fb2 : _GEN_2506; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2508 = 5'h15 == _T_280[4:0] ? 32'h3f800000 : _GEN_2507; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2509 = 5'h16 == _T_280[4:0] ? 32'hbd6e2940 : _GEN_2508; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2510 = 5'h17 == _T_280[4:0] ? 32'hbf7e44de : _GEN_2509; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2511 = 5'h18 == _T_280[4:0] ? 32'h3f800000 : _GEN_2510; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2512 = 5'h19 == _T_280[4:0] ? 32'hbe92d7dc : _GEN_2511; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2518 = 5'h4 == _T_280[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2519 = 5'h5 == _T_280[4:0] ? 32'hbee5c900 : _GEN_2518; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2520 = 5'h6 == _T_280[4:0] ? 32'h80800000 : _GEN_2519; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2521 = 5'h7 == _T_280[4:0] ? 32'hbee5c900 : _GEN_2520; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2522 = 5'h8 == _T_280[4:0] ? 32'hbf4d57f2 : _GEN_2521; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2523 = 5'h9 == _T_280[4:0] ? 32'h80800000 : _GEN_2522; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2524 = 5'ha == _T_280[4:0] ? 32'hbf248dba : _GEN_2523; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2525 = 5'hb == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2524; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2526 = 5'hc == _T_280[4:0] ? 32'h80800000 : _GEN_2525; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2527 = 5'hd == _T_280[4:0] ? 32'hbf4d57f2 : _GEN_2526; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2528 = 5'he == _T_280[4:0] ? 32'hbf753ecc : _GEN_2527; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2529 = 5'hf == _T_280[4:0] ? 32'h80800000 : _GEN_2528; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2530 = 5'h10 == _T_280[4:0] ? 32'hbf6b1034 : _GEN_2529; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2531 = 5'h11 == _T_280[4:0] ? 32'hbf3a3528 : _GEN_2530; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2532 = 5'h12 == _T_280[4:0] ? 32'h80800000 : _GEN_2531; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2533 = 5'h13 == _T_280[4:0] ? 32'hbf7c1c5c : _GEN_2532; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2534 = 5'h14 == _T_280[4:0] ? 32'hbeaf1d40 : _GEN_2533; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2535 = 5'h15 == _T_280[4:0] ? 32'h80800000 : _GEN_2534; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2536 = 5'h16 == _T_280[4:0] ? 32'hbf7f911e : _GEN_2535; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2537 = 5'h17 == _T_280[4:0] ? 32'h3dedc210 : _GEN_2536; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2538 = 5'h18 == _T_280[4:0] ? 32'h80800000 : _GEN_2537; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2539 = 5'h19 == _T_280[4:0] ? 32'hbf753ecc : _GEN_2538; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2542 = 5'h1 == _T_280[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2543 = 5'h2 == _T_280[4:0] ? io_in_2_Im : _GEN_2542; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2544 = 5'h3 == _T_280[4:0] ? io_in_3_Im : _GEN_2543; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2545 = 5'h4 == _T_280[4:0] ? io_in_4_Im : _GEN_2544; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2546 = 5'h5 == _T_280[4:0] ? io_in_5_Im : _GEN_2545; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2547 = 5'h6 == _T_280[4:0] ? io_in_6_Im : _GEN_2546; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2548 = 5'h7 == _T_280[4:0] ? io_in_7_Im : _GEN_2547; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2549 = 5'h8 == _T_280[4:0] ? io_in_8_Im : _GEN_2548; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2550 = 5'h9 == _T_280[4:0] ? io_in_9_Im : _GEN_2549; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2551 = 5'ha == _T_280[4:0] ? io_in_10_Im : _GEN_2550; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2552 = 5'hb == _T_280[4:0] ? io_in_11_Im : _GEN_2551; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2553 = 5'hc == _T_280[4:0] ? io_in_12_Im : _GEN_2552; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2554 = 5'hd == _T_280[4:0] ? io_in_13_Im : _GEN_2553; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2555 = 5'he == _T_280[4:0] ? io_in_14_Im : _GEN_2554; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2556 = 5'hf == _T_280[4:0] ? io_in_15_Im : _GEN_2555; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2557 = 5'h10 == _T_280[4:0] ? io_in_16_Im : _GEN_2556; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2558 = 5'h11 == _T_280[4:0] ? io_in_17_Im : _GEN_2557; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2559 = 5'h12 == _T_280[4:0] ? io_in_18_Im : _GEN_2558; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2560 = 5'h13 == _T_280[4:0] ? io_in_19_Im : _GEN_2559; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2561 = 5'h14 == _T_280[4:0] ? io_in_20_Im : _GEN_2560; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2562 = 5'h15 == _T_280[4:0] ? io_in_21_Im : _GEN_2561; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2563 = 5'h16 == _T_280[4:0] ? io_in_22_Im : _GEN_2562; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2564 = 5'h17 == _T_280[4:0] ? io_in_23_Im : _GEN_2563; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2565 = 5'h18 == _T_280[4:0] ? io_in_24_Im : _GEN_2564; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2566 = 5'h19 == _T_280[4:0] ? io_in_25_Im : _GEN_2565; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2569 = 5'h1 == _T_280[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2570 = 5'h2 == _T_280[4:0] ? io_in_2_Re : _GEN_2569; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2571 = 5'h3 == _T_280[4:0] ? io_in_3_Re : _GEN_2570; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2572 = 5'h4 == _T_280[4:0] ? io_in_4_Re : _GEN_2571; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2573 = 5'h5 == _T_280[4:0] ? io_in_5_Re : _GEN_2572; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2574 = 5'h6 == _T_280[4:0] ? io_in_6_Re : _GEN_2573; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2575 = 5'h7 == _T_280[4:0] ? io_in_7_Re : _GEN_2574; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2576 = 5'h8 == _T_280[4:0] ? io_in_8_Re : _GEN_2575; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2577 = 5'h9 == _T_280[4:0] ? io_in_9_Re : _GEN_2576; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2578 = 5'ha == _T_280[4:0] ? io_in_10_Re : _GEN_2577; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2579 = 5'hb == _T_280[4:0] ? io_in_11_Re : _GEN_2578; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2580 = 5'hc == _T_280[4:0] ? io_in_12_Re : _GEN_2579; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2581 = 5'hd == _T_280[4:0] ? io_in_13_Re : _GEN_2580; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2582 = 5'he == _T_280[4:0] ? io_in_14_Re : _GEN_2581; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2583 = 5'hf == _T_280[4:0] ? io_in_15_Re : _GEN_2582; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2584 = 5'h10 == _T_280[4:0] ? io_in_16_Re : _GEN_2583; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2585 = 5'h11 == _T_280[4:0] ? io_in_17_Re : _GEN_2584; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2586 = 5'h12 == _T_280[4:0] ? io_in_18_Re : _GEN_2585; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2587 = 5'h13 == _T_280[4:0] ? io_in_19_Re : _GEN_2586; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2588 = 5'h14 == _T_280[4:0] ? io_in_20_Re : _GEN_2587; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2589 = 5'h15 == _T_280[4:0] ? io_in_21_Re : _GEN_2588; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2590 = 5'h16 == _T_280[4:0] ? io_in_22_Re : _GEN_2589; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2591 = 5'h17 == _T_280[4:0] ? io_in_23_Re : _GEN_2590; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2592 = 5'h18 == _T_280[4:0] ? io_in_24_Re : _GEN_2591; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2593 = 5'h19 == _T_280[4:0] ? io_in_25_Re : _GEN_2592; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_292 = _T_2 + 37'h18; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2599 = 5'h4 == _T_292[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2600 = 5'h5 == _T_292[4:0] ? 32'h3f64c51a : _GEN_2599; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2601 = 5'h6 == _T_292[4:0] ? 32'h3f800000 : _GEN_2600; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2602 = 5'h7 == _T_292[4:0] ? 32'h3f64c51a : _GEN_2601; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2603 = 5'h8 == _T_292[4:0] ? 32'h3f18df62 : _GEN_2602; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2604 = 5'h9 == _T_292[4:0] ? 32'h3f800000 : _GEN_2603; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2605 = 5'ha == _T_292[4:0] ? 32'h3f441b7c : _GEN_2604; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2606 = 5'hb == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2605; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2607 = 5'hc == _T_292[4:0] ? 32'h3f800000 : _GEN_2606; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2608 = 5'hd == _T_292[4:0] ? 32'h3f18df62 : _GEN_2607; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2609 = 5'he == _T_292[4:0] ? 32'hbe92d7dc : _GEN_2608; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2610 = 5'hf == _T_292[4:0] ? 32'h3f800000 : _GEN_2609; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2611 = 5'h10 == _T_292[4:0] ? 32'h3ecacaf4 : _GEN_2610; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2612 = 5'h11 == _T_292[4:0] ? 32'hbf2fad88 : _GEN_2611; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2613 = 5'h12 == _T_292[4:0] ? 32'h3f800000 : _GEN_2612; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2614 = 5'h13 == _T_292[4:0] ? 32'h3e31d0d0 : _GEN_2613; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2615 = 5'h14 == _T_292[4:0] ? 32'hbf708fb2 : _GEN_2614; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2616 = 5'h15 == _T_292[4:0] ? 32'h3f800000 : _GEN_2615; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2617 = 5'h16 == _T_292[4:0] ? 32'hbd6e2940 : _GEN_2616; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2618 = 5'h17 == _T_292[4:0] ? 32'hbf7e44de : _GEN_2617; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2619 = 5'h18 == _T_292[4:0] ? 32'h3f800000 : _GEN_2618; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2620 = 5'h19 == _T_292[4:0] ? 32'hbe92d7dc : _GEN_2619; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2626 = 5'h4 == _T_292[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2627 = 5'h5 == _T_292[4:0] ? 32'hbee5c900 : _GEN_2626; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2628 = 5'h6 == _T_292[4:0] ? 32'h80800000 : _GEN_2627; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2629 = 5'h7 == _T_292[4:0] ? 32'hbee5c900 : _GEN_2628; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2630 = 5'h8 == _T_292[4:0] ? 32'hbf4d57f2 : _GEN_2629; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2631 = 5'h9 == _T_292[4:0] ? 32'h80800000 : _GEN_2630; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2632 = 5'ha == _T_292[4:0] ? 32'hbf248dba : _GEN_2631; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2633 = 5'hb == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2632; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2634 = 5'hc == _T_292[4:0] ? 32'h80800000 : _GEN_2633; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2635 = 5'hd == _T_292[4:0] ? 32'hbf4d57f2 : _GEN_2634; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2636 = 5'he == _T_292[4:0] ? 32'hbf753ecc : _GEN_2635; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2637 = 5'hf == _T_292[4:0] ? 32'h80800000 : _GEN_2636; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2638 = 5'h10 == _T_292[4:0] ? 32'hbf6b1034 : _GEN_2637; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2639 = 5'h11 == _T_292[4:0] ? 32'hbf3a3528 : _GEN_2638; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2640 = 5'h12 == _T_292[4:0] ? 32'h80800000 : _GEN_2639; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2641 = 5'h13 == _T_292[4:0] ? 32'hbf7c1c5c : _GEN_2640; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2642 = 5'h14 == _T_292[4:0] ? 32'hbeaf1d40 : _GEN_2641; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2643 = 5'h15 == _T_292[4:0] ? 32'h80800000 : _GEN_2642; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2644 = 5'h16 == _T_292[4:0] ? 32'hbf7f911e : _GEN_2643; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2645 = 5'h17 == _T_292[4:0] ? 32'h3dedc210 : _GEN_2644; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2646 = 5'h18 == _T_292[4:0] ? 32'h80800000 : _GEN_2645; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2647 = 5'h19 == _T_292[4:0] ? 32'hbf753ecc : _GEN_2646; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2650 = 5'h1 == _T_292[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2651 = 5'h2 == _T_292[4:0] ? io_in_2_Im : _GEN_2650; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2652 = 5'h3 == _T_292[4:0] ? io_in_3_Im : _GEN_2651; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2653 = 5'h4 == _T_292[4:0] ? io_in_4_Im : _GEN_2652; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2654 = 5'h5 == _T_292[4:0] ? io_in_5_Im : _GEN_2653; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2655 = 5'h6 == _T_292[4:0] ? io_in_6_Im : _GEN_2654; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2656 = 5'h7 == _T_292[4:0] ? io_in_7_Im : _GEN_2655; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2657 = 5'h8 == _T_292[4:0] ? io_in_8_Im : _GEN_2656; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2658 = 5'h9 == _T_292[4:0] ? io_in_9_Im : _GEN_2657; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2659 = 5'ha == _T_292[4:0] ? io_in_10_Im : _GEN_2658; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2660 = 5'hb == _T_292[4:0] ? io_in_11_Im : _GEN_2659; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2661 = 5'hc == _T_292[4:0] ? io_in_12_Im : _GEN_2660; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2662 = 5'hd == _T_292[4:0] ? io_in_13_Im : _GEN_2661; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2663 = 5'he == _T_292[4:0] ? io_in_14_Im : _GEN_2662; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2664 = 5'hf == _T_292[4:0] ? io_in_15_Im : _GEN_2663; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2665 = 5'h10 == _T_292[4:0] ? io_in_16_Im : _GEN_2664; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2666 = 5'h11 == _T_292[4:0] ? io_in_17_Im : _GEN_2665; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2667 = 5'h12 == _T_292[4:0] ? io_in_18_Im : _GEN_2666; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2668 = 5'h13 == _T_292[4:0] ? io_in_19_Im : _GEN_2667; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2669 = 5'h14 == _T_292[4:0] ? io_in_20_Im : _GEN_2668; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2670 = 5'h15 == _T_292[4:0] ? io_in_21_Im : _GEN_2669; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2671 = 5'h16 == _T_292[4:0] ? io_in_22_Im : _GEN_2670; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2672 = 5'h17 == _T_292[4:0] ? io_in_23_Im : _GEN_2671; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2673 = 5'h18 == _T_292[4:0] ? io_in_24_Im : _GEN_2672; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2674 = 5'h19 == _T_292[4:0] ? io_in_25_Im : _GEN_2673; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2677 = 5'h1 == _T_292[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2678 = 5'h2 == _T_292[4:0] ? io_in_2_Re : _GEN_2677; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2679 = 5'h3 == _T_292[4:0] ? io_in_3_Re : _GEN_2678; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2680 = 5'h4 == _T_292[4:0] ? io_in_4_Re : _GEN_2679; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2681 = 5'h5 == _T_292[4:0] ? io_in_5_Re : _GEN_2680; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2682 = 5'h6 == _T_292[4:0] ? io_in_6_Re : _GEN_2681; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2683 = 5'h7 == _T_292[4:0] ? io_in_7_Re : _GEN_2682; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2684 = 5'h8 == _T_292[4:0] ? io_in_8_Re : _GEN_2683; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2685 = 5'h9 == _T_292[4:0] ? io_in_9_Re : _GEN_2684; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2686 = 5'ha == _T_292[4:0] ? io_in_10_Re : _GEN_2685; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2687 = 5'hb == _T_292[4:0] ? io_in_11_Re : _GEN_2686; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2688 = 5'hc == _T_292[4:0] ? io_in_12_Re : _GEN_2687; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2689 = 5'hd == _T_292[4:0] ? io_in_13_Re : _GEN_2688; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2690 = 5'he == _T_292[4:0] ? io_in_14_Re : _GEN_2689; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2691 = 5'hf == _T_292[4:0] ? io_in_15_Re : _GEN_2690; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2692 = 5'h10 == _T_292[4:0] ? io_in_16_Re : _GEN_2691; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2693 = 5'h11 == _T_292[4:0] ? io_in_17_Re : _GEN_2692; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2694 = 5'h12 == _T_292[4:0] ? io_in_18_Re : _GEN_2693; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2695 = 5'h13 == _T_292[4:0] ? io_in_19_Re : _GEN_2694; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2696 = 5'h14 == _T_292[4:0] ? io_in_20_Re : _GEN_2695; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2697 = 5'h15 == _T_292[4:0] ? io_in_21_Re : _GEN_2696; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2698 = 5'h16 == _T_292[4:0] ? io_in_22_Re : _GEN_2697; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2699 = 5'h17 == _T_292[4:0] ? io_in_23_Re : _GEN_2698; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2700 = 5'h18 == _T_292[4:0] ? io_in_24_Re : _GEN_2699; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2701 = 5'h19 == _T_292[4:0] ? io_in_25_Re : _GEN_2700; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_304 = _T_2 + 37'h19; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2707 = 5'h4 == _T_304[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2708 = 5'h5 == _T_304[4:0] ? 32'h3f64c51a : _GEN_2707; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2709 = 5'h6 == _T_304[4:0] ? 32'h3f800000 : _GEN_2708; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2710 = 5'h7 == _T_304[4:0] ? 32'h3f64c51a : _GEN_2709; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2711 = 5'h8 == _T_304[4:0] ? 32'h3f18df62 : _GEN_2710; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2712 = 5'h9 == _T_304[4:0] ? 32'h3f800000 : _GEN_2711; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2713 = 5'ha == _T_304[4:0] ? 32'h3f441b7c : _GEN_2712; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2714 = 5'hb == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2713; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2715 = 5'hc == _T_304[4:0] ? 32'h3f800000 : _GEN_2714; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2716 = 5'hd == _T_304[4:0] ? 32'h3f18df62 : _GEN_2715; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2717 = 5'he == _T_304[4:0] ? 32'hbe92d7dc : _GEN_2716; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2718 = 5'hf == _T_304[4:0] ? 32'h3f800000 : _GEN_2717; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2719 = 5'h10 == _T_304[4:0] ? 32'h3ecacaf4 : _GEN_2718; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2720 = 5'h11 == _T_304[4:0] ? 32'hbf2fad88 : _GEN_2719; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2721 = 5'h12 == _T_304[4:0] ? 32'h3f800000 : _GEN_2720; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2722 = 5'h13 == _T_304[4:0] ? 32'h3e31d0d0 : _GEN_2721; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2723 = 5'h14 == _T_304[4:0] ? 32'hbf708fb2 : _GEN_2722; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2724 = 5'h15 == _T_304[4:0] ? 32'h3f800000 : _GEN_2723; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2725 = 5'h16 == _T_304[4:0] ? 32'hbd6e2940 : _GEN_2724; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2726 = 5'h17 == _T_304[4:0] ? 32'hbf7e44de : _GEN_2725; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2727 = 5'h18 == _T_304[4:0] ? 32'h3f800000 : _GEN_2726; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2728 = 5'h19 == _T_304[4:0] ? 32'hbe92d7dc : _GEN_2727; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2734 = 5'h4 == _T_304[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2735 = 5'h5 == _T_304[4:0] ? 32'hbee5c900 : _GEN_2734; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2736 = 5'h6 == _T_304[4:0] ? 32'h80800000 : _GEN_2735; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2737 = 5'h7 == _T_304[4:0] ? 32'hbee5c900 : _GEN_2736; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2738 = 5'h8 == _T_304[4:0] ? 32'hbf4d57f2 : _GEN_2737; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2739 = 5'h9 == _T_304[4:0] ? 32'h80800000 : _GEN_2738; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2740 = 5'ha == _T_304[4:0] ? 32'hbf248dba : _GEN_2739; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2741 = 5'hb == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2740; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2742 = 5'hc == _T_304[4:0] ? 32'h80800000 : _GEN_2741; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2743 = 5'hd == _T_304[4:0] ? 32'hbf4d57f2 : _GEN_2742; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2744 = 5'he == _T_304[4:0] ? 32'hbf753ecc : _GEN_2743; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2745 = 5'hf == _T_304[4:0] ? 32'h80800000 : _GEN_2744; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2746 = 5'h10 == _T_304[4:0] ? 32'hbf6b1034 : _GEN_2745; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2747 = 5'h11 == _T_304[4:0] ? 32'hbf3a3528 : _GEN_2746; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2748 = 5'h12 == _T_304[4:0] ? 32'h80800000 : _GEN_2747; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2749 = 5'h13 == _T_304[4:0] ? 32'hbf7c1c5c : _GEN_2748; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2750 = 5'h14 == _T_304[4:0] ? 32'hbeaf1d40 : _GEN_2749; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2751 = 5'h15 == _T_304[4:0] ? 32'h80800000 : _GEN_2750; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2752 = 5'h16 == _T_304[4:0] ? 32'hbf7f911e : _GEN_2751; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2753 = 5'h17 == _T_304[4:0] ? 32'h3dedc210 : _GEN_2752; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2754 = 5'h18 == _T_304[4:0] ? 32'h80800000 : _GEN_2753; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2755 = 5'h19 == _T_304[4:0] ? 32'hbf753ecc : _GEN_2754; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2758 = 5'h1 == _T_304[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2759 = 5'h2 == _T_304[4:0] ? io_in_2_Im : _GEN_2758; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2760 = 5'h3 == _T_304[4:0] ? io_in_3_Im : _GEN_2759; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2761 = 5'h4 == _T_304[4:0] ? io_in_4_Im : _GEN_2760; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2762 = 5'h5 == _T_304[4:0] ? io_in_5_Im : _GEN_2761; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2763 = 5'h6 == _T_304[4:0] ? io_in_6_Im : _GEN_2762; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2764 = 5'h7 == _T_304[4:0] ? io_in_7_Im : _GEN_2763; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2765 = 5'h8 == _T_304[4:0] ? io_in_8_Im : _GEN_2764; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2766 = 5'h9 == _T_304[4:0] ? io_in_9_Im : _GEN_2765; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2767 = 5'ha == _T_304[4:0] ? io_in_10_Im : _GEN_2766; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2768 = 5'hb == _T_304[4:0] ? io_in_11_Im : _GEN_2767; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2769 = 5'hc == _T_304[4:0] ? io_in_12_Im : _GEN_2768; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2770 = 5'hd == _T_304[4:0] ? io_in_13_Im : _GEN_2769; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2771 = 5'he == _T_304[4:0] ? io_in_14_Im : _GEN_2770; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2772 = 5'hf == _T_304[4:0] ? io_in_15_Im : _GEN_2771; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2773 = 5'h10 == _T_304[4:0] ? io_in_16_Im : _GEN_2772; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2774 = 5'h11 == _T_304[4:0] ? io_in_17_Im : _GEN_2773; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2775 = 5'h12 == _T_304[4:0] ? io_in_18_Im : _GEN_2774; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2776 = 5'h13 == _T_304[4:0] ? io_in_19_Im : _GEN_2775; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2777 = 5'h14 == _T_304[4:0] ? io_in_20_Im : _GEN_2776; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2778 = 5'h15 == _T_304[4:0] ? io_in_21_Im : _GEN_2777; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2779 = 5'h16 == _T_304[4:0] ? io_in_22_Im : _GEN_2778; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2780 = 5'h17 == _T_304[4:0] ? io_in_23_Im : _GEN_2779; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2781 = 5'h18 == _T_304[4:0] ? io_in_24_Im : _GEN_2780; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2782 = 5'h19 == _T_304[4:0] ? io_in_25_Im : _GEN_2781; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2785 = 5'h1 == _T_304[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2786 = 5'h2 == _T_304[4:0] ? io_in_2_Re : _GEN_2785; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2787 = 5'h3 == _T_304[4:0] ? io_in_3_Re : _GEN_2786; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2788 = 5'h4 == _T_304[4:0] ? io_in_4_Re : _GEN_2787; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2789 = 5'h5 == _T_304[4:0] ? io_in_5_Re : _GEN_2788; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2790 = 5'h6 == _T_304[4:0] ? io_in_6_Re : _GEN_2789; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2791 = 5'h7 == _T_304[4:0] ? io_in_7_Re : _GEN_2790; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2792 = 5'h8 == _T_304[4:0] ? io_in_8_Re : _GEN_2791; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2793 = 5'h9 == _T_304[4:0] ? io_in_9_Re : _GEN_2792; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2794 = 5'ha == _T_304[4:0] ? io_in_10_Re : _GEN_2793; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2795 = 5'hb == _T_304[4:0] ? io_in_11_Re : _GEN_2794; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2796 = 5'hc == _T_304[4:0] ? io_in_12_Re : _GEN_2795; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2797 = 5'hd == _T_304[4:0] ? io_in_13_Re : _GEN_2796; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2798 = 5'he == _T_304[4:0] ? io_in_14_Re : _GEN_2797; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2799 = 5'hf == _T_304[4:0] ? io_in_15_Re : _GEN_2798; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2800 = 5'h10 == _T_304[4:0] ? io_in_16_Re : _GEN_2799; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2801 = 5'h11 == _T_304[4:0] ? io_in_17_Re : _GEN_2800; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2802 = 5'h12 == _T_304[4:0] ? io_in_18_Re : _GEN_2801; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2803 = 5'h13 == _T_304[4:0] ? io_in_19_Re : _GEN_2802; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2804 = 5'h14 == _T_304[4:0] ? io_in_20_Re : _GEN_2803; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2805 = 5'h15 == _T_304[4:0] ? io_in_21_Re : _GEN_2804; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2806 = 5'h16 == _T_304[4:0] ? io_in_22_Re : _GEN_2805; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2807 = 5'h17 == _T_304[4:0] ? io_in_23_Re : _GEN_2806; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2808 = 5'h18 == _T_304[4:0] ? io_in_24_Re : _GEN_2807; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2809 = 5'h19 == _T_304[4:0] ? io_in_25_Re : _GEN_2808; // @[FFTDesigns.scala 543:{23,23}]
  wire [36:0] _T_316 = _T_2 + 37'h1a; // @[FFTDesigns.scala 541:64]
  wire [31:0] _GEN_2815 = 5'h4 == _T_316[4:0] ? 32'h3f791976 : 32'h3f800000; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2816 = 5'h5 == _T_316[4:0] ? 32'h3f64c51a : _GEN_2815; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2817 = 5'h6 == _T_316[4:0] ? 32'h3f800000 : _GEN_2816; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2818 = 5'h7 == _T_316[4:0] ? 32'h3f64c51a : _GEN_2817; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2819 = 5'h8 == _T_316[4:0] ? 32'h3f18df62 : _GEN_2818; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2820 = 5'h9 == _T_316[4:0] ? 32'h3f800000 : _GEN_2819; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2821 = 5'ha == _T_316[4:0] ? 32'h3f441b7c : _GEN_2820; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2822 = 5'hb == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2821; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2823 = 5'hc == _T_316[4:0] ? 32'h3f800000 : _GEN_2822; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2824 = 5'hd == _T_316[4:0] ? 32'h3f18df62 : _GEN_2823; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2825 = 5'he == _T_316[4:0] ? 32'hbe92d7dc : _GEN_2824; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2826 = 5'hf == _T_316[4:0] ? 32'h3f800000 : _GEN_2825; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2827 = 5'h10 == _T_316[4:0] ? 32'h3ecacaf4 : _GEN_2826; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2828 = 5'h11 == _T_316[4:0] ? 32'hbf2fad88 : _GEN_2827; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2829 = 5'h12 == _T_316[4:0] ? 32'h3f800000 : _GEN_2828; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2830 = 5'h13 == _T_316[4:0] ? 32'h3e31d0d0 : _GEN_2829; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2831 = 5'h14 == _T_316[4:0] ? 32'hbf708fb2 : _GEN_2830; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2832 = 5'h15 == _T_316[4:0] ? 32'h3f800000 : _GEN_2831; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2833 = 5'h16 == _T_316[4:0] ? 32'hbd6e2940 : _GEN_2832; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2834 = 5'h17 == _T_316[4:0] ? 32'hbf7e44de : _GEN_2833; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2835 = 5'h18 == _T_316[4:0] ? 32'h3f800000 : _GEN_2834; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2836 = 5'h19 == _T_316[4:0] ? 32'hbe92d7dc : _GEN_2835; // @[FFTDesigns.scala 541:{26,26}]
  wire [31:0] _GEN_2842 = 5'h4 == _T_316[4:0] ? 32'hbe6c2690 : 32'h80800000; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2843 = 5'h5 == _T_316[4:0] ? 32'hbee5c900 : _GEN_2842; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2844 = 5'h6 == _T_316[4:0] ? 32'h80800000 : _GEN_2843; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2845 = 5'h7 == _T_316[4:0] ? 32'hbee5c900 : _GEN_2844; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2846 = 5'h8 == _T_316[4:0] ? 32'hbf4d57f2 : _GEN_2845; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2847 = 5'h9 == _T_316[4:0] ? 32'h80800000 : _GEN_2846; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2848 = 5'ha == _T_316[4:0] ? 32'hbf248dba : _GEN_2847; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2849 = 5'hb == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2848; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2850 = 5'hc == _T_316[4:0] ? 32'h80800000 : _GEN_2849; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2851 = 5'hd == _T_316[4:0] ? 32'hbf4d57f2 : _GEN_2850; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2852 = 5'he == _T_316[4:0] ? 32'hbf753ecc : _GEN_2851; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2853 = 5'hf == _T_316[4:0] ? 32'h80800000 : _GEN_2852; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2854 = 5'h10 == _T_316[4:0] ? 32'hbf6b1034 : _GEN_2853; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2855 = 5'h11 == _T_316[4:0] ? 32'hbf3a3528 : _GEN_2854; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2856 = 5'h12 == _T_316[4:0] ? 32'h80800000 : _GEN_2855; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2857 = 5'h13 == _T_316[4:0] ? 32'hbf7c1c5c : _GEN_2856; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2858 = 5'h14 == _T_316[4:0] ? 32'hbeaf1d40 : _GEN_2857; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2859 = 5'h15 == _T_316[4:0] ? 32'h80800000 : _GEN_2858; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2860 = 5'h16 == _T_316[4:0] ? 32'hbf7f911e : _GEN_2859; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2861 = 5'h17 == _T_316[4:0] ? 32'h3dedc210 : _GEN_2860; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2862 = 5'h18 == _T_316[4:0] ? 32'h80800000 : _GEN_2861; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2863 = 5'h19 == _T_316[4:0] ? 32'hbf753ecc : _GEN_2862; // @[FFTDesigns.scala 542:{26,26}]
  wire [31:0] _GEN_2866 = 5'h1 == _T_316[4:0] ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2867 = 5'h2 == _T_316[4:0] ? io_in_2_Im : _GEN_2866; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2868 = 5'h3 == _T_316[4:0] ? io_in_3_Im : _GEN_2867; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2869 = 5'h4 == _T_316[4:0] ? io_in_4_Im : _GEN_2868; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2870 = 5'h5 == _T_316[4:0] ? io_in_5_Im : _GEN_2869; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2871 = 5'h6 == _T_316[4:0] ? io_in_6_Im : _GEN_2870; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2872 = 5'h7 == _T_316[4:0] ? io_in_7_Im : _GEN_2871; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2873 = 5'h8 == _T_316[4:0] ? io_in_8_Im : _GEN_2872; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2874 = 5'h9 == _T_316[4:0] ? io_in_9_Im : _GEN_2873; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2875 = 5'ha == _T_316[4:0] ? io_in_10_Im : _GEN_2874; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2876 = 5'hb == _T_316[4:0] ? io_in_11_Im : _GEN_2875; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2877 = 5'hc == _T_316[4:0] ? io_in_12_Im : _GEN_2876; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2878 = 5'hd == _T_316[4:0] ? io_in_13_Im : _GEN_2877; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2879 = 5'he == _T_316[4:0] ? io_in_14_Im : _GEN_2878; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2880 = 5'hf == _T_316[4:0] ? io_in_15_Im : _GEN_2879; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2881 = 5'h10 == _T_316[4:0] ? io_in_16_Im : _GEN_2880; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2882 = 5'h11 == _T_316[4:0] ? io_in_17_Im : _GEN_2881; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2883 = 5'h12 == _T_316[4:0] ? io_in_18_Im : _GEN_2882; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2884 = 5'h13 == _T_316[4:0] ? io_in_19_Im : _GEN_2883; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2885 = 5'h14 == _T_316[4:0] ? io_in_20_Im : _GEN_2884; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2886 = 5'h15 == _T_316[4:0] ? io_in_21_Im : _GEN_2885; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2887 = 5'h16 == _T_316[4:0] ? io_in_22_Im : _GEN_2886; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2888 = 5'h17 == _T_316[4:0] ? io_in_23_Im : _GEN_2887; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2889 = 5'h18 == _T_316[4:0] ? io_in_24_Im : _GEN_2888; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2890 = 5'h19 == _T_316[4:0] ? io_in_25_Im : _GEN_2889; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2893 = 5'h1 == _T_316[4:0] ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2894 = 5'h2 == _T_316[4:0] ? io_in_2_Re : _GEN_2893; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2895 = 5'h3 == _T_316[4:0] ? io_in_3_Re : _GEN_2894; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2896 = 5'h4 == _T_316[4:0] ? io_in_4_Re : _GEN_2895; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2897 = 5'h5 == _T_316[4:0] ? io_in_5_Re : _GEN_2896; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2898 = 5'h6 == _T_316[4:0] ? io_in_6_Re : _GEN_2897; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2899 = 5'h7 == _T_316[4:0] ? io_in_7_Re : _GEN_2898; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2900 = 5'h8 == _T_316[4:0] ? io_in_8_Re : _GEN_2899; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2901 = 5'h9 == _T_316[4:0] ? io_in_9_Re : _GEN_2900; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2902 = 5'ha == _T_316[4:0] ? io_in_10_Re : _GEN_2901; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2903 = 5'hb == _T_316[4:0] ? io_in_11_Re : _GEN_2902; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2904 = 5'hc == _T_316[4:0] ? io_in_12_Re : _GEN_2903; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2905 = 5'hd == _T_316[4:0] ? io_in_13_Re : _GEN_2904; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2906 = 5'he == _T_316[4:0] ? io_in_14_Re : _GEN_2905; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2907 = 5'hf == _T_316[4:0] ? io_in_15_Re : _GEN_2906; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2908 = 5'h10 == _T_316[4:0] ? io_in_16_Re : _GEN_2907; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2909 = 5'h11 == _T_316[4:0] ? io_in_17_Re : _GEN_2908; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2910 = 5'h12 == _T_316[4:0] ? io_in_18_Re : _GEN_2909; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2911 = 5'h13 == _T_316[4:0] ? io_in_19_Re : _GEN_2910; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2912 = 5'h14 == _T_316[4:0] ? io_in_20_Re : _GEN_2911; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2913 = 5'h15 == _T_316[4:0] ? io_in_21_Re : _GEN_2912; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2914 = 5'h16 == _T_316[4:0] ? io_in_22_Re : _GEN_2913; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2915 = 5'h17 == _T_316[4:0] ? io_in_23_Re : _GEN_2914; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2916 = 5'h18 == _T_316[4:0] ? io_in_24_Re : _GEN_2915; // @[FFTDesigns.scala 543:{23,23}]
  wire [31:0] _GEN_2917 = 5'h19 == _T_316[4:0] ? io_in_25_Re : _GEN_2916; // @[FFTDesigns.scala 543:{23,23}]
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_clock),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_1_clock),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_2_clock),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_3_clock),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_4_clock),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_5_clock),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_6_clock),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_7_clock),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_8_clock),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_9_clock),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_10_clock),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_11_clock),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_12 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_12_clock),
    .io_in_a_Re(FPComplexMult_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_12_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_13 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_13_clock),
    .io_in_a_Re(FPComplexMult_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_13_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_14 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_14_clock),
    .io_in_a_Re(FPComplexMult_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_14_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_15 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_15_clock),
    .io_in_a_Re(FPComplexMult_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_15_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_16 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_16_clock),
    .io_in_a_Re(FPComplexMult_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_16_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_16_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_16_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_16_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_17 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_17_clock),
    .io_in_a_Re(FPComplexMult_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_17_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_17_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_17_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_17_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_18 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_18_clock),
    .io_in_a_Re(FPComplexMult_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_18_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_18_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_18_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_18_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_19 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_19_clock),
    .io_in_a_Re(FPComplexMult_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_19_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_19_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_19_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_19_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_20 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_20_clock),
    .io_in_a_Re(FPComplexMult_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_20_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_20_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_20_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_20_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_21 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_21_clock),
    .io_in_a_Re(FPComplexMult_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_21_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_21_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_21_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_21_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_22 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_22_clock),
    .io_in_a_Re(FPComplexMult_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_22_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_22_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_22_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_22_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_23 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_23_clock),
    .io_in_a_Re(FPComplexMult_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_23_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_23_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_23_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_23_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_24 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_24_clock),
    .io_in_a_Re(FPComplexMult_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_24_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_24_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_24_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_24_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_25 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_25_clock),
    .io_in_a_Re(FPComplexMult_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_25_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_25_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_25_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_25_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_26 ( // @[FFTDesigns.scala 524:26]
    .clock(FPComplexMult_26_clock),
    .io_in_a_Re(FPComplexMult_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_26_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_26_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_26_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_26_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_12_Re = FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_12_Im = FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_13_Re = FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_13_Im = FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_14_Re = FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_14_Im = FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_15_Re = FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_15_Im = FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_16_Re = FPComplexMult_16_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_16_Im = FPComplexMult_16_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_17_Re = FPComplexMult_17_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_17_Im = FPComplexMult_17_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_18_Re = FPComplexMult_18_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_18_Im = FPComplexMult_18_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_19_Re = FPComplexMult_19_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_19_Im = FPComplexMult_19_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_20_Re = FPComplexMult_20_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_20_Im = FPComplexMult_20_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_21_Re = FPComplexMult_21_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_21_Im = FPComplexMult_21_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_22_Re = FPComplexMult_22_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_22_Im = FPComplexMult_22_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_23_Re = FPComplexMult_23_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_23_Im = FPComplexMult_23_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_24_Re = FPComplexMult_24_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_24_Im = FPComplexMult_24_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_25_Re = FPComplexMult_25_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_25_Im = FPComplexMult_25_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign io_out_26_Re = FPComplexMult_26_io_out_s_Re; // @[FFTDesigns.scala 544:17]
  assign io_out_26_Im = FPComplexMult_26_io_out_s_Im; // @[FFTDesigns.scala 544:17]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_io_in_a_Re = 5'h1a == _T_3[4:0] ? 32'hbf55e286 : _GEN_28; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_io_in_a_Im = 5'h1a == _T_3[4:0] ? 32'h3f0cac9e : _GEN_55; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_io_in_b_Re = 5'h1a == _T_3[4:0] ? io_in_26_Re : _GEN_109; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_io_in_b_Im = 5'h1a == _T_3[4:0] ? io_in_26_Im : _GEN_82; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_io_in_a_Re = 5'h1a == _T_16[4:0] ? 32'hbf55e286 : _GEN_136; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_1_io_in_a_Im = 5'h1a == _T_16[4:0] ? 32'h3f0cac9e : _GEN_163; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_1_io_in_b_Re = 5'h1a == _T_16[4:0] ? io_in_26_Re : _GEN_217; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_1_io_in_b_Im = 5'h1a == _T_16[4:0] ? io_in_26_Im : _GEN_190; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_io_in_a_Re = 5'h1a == _T_28[4:0] ? 32'hbf55e286 : _GEN_244; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_2_io_in_a_Im = 5'h1a == _T_28[4:0] ? 32'h3f0cac9e : _GEN_271; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_2_io_in_b_Re = 5'h1a == _T_28[4:0] ? io_in_26_Re : _GEN_325; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_2_io_in_b_Im = 5'h1a == _T_28[4:0] ? io_in_26_Im : _GEN_298; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_io_in_a_Re = 5'h1a == _T_40[4:0] ? 32'hbf55e286 : _GEN_352; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_3_io_in_a_Im = 5'h1a == _T_40[4:0] ? 32'h3f0cac9e : _GEN_379; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_3_io_in_b_Re = 5'h1a == _T_40[4:0] ? io_in_26_Re : _GEN_433; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_3_io_in_b_Im = 5'h1a == _T_40[4:0] ? io_in_26_Im : _GEN_406; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_io_in_a_Re = 5'h1a == _T_52[4:0] ? 32'hbf55e286 : _GEN_460; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_4_io_in_a_Im = 5'h1a == _T_52[4:0] ? 32'h3f0cac9e : _GEN_487; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_4_io_in_b_Re = 5'h1a == _T_52[4:0] ? io_in_26_Re : _GEN_541; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_4_io_in_b_Im = 5'h1a == _T_52[4:0] ? io_in_26_Im : _GEN_514; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_io_in_a_Re = 5'h1a == _T_64[4:0] ? 32'hbf55e286 : _GEN_568; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_5_io_in_a_Im = 5'h1a == _T_64[4:0] ? 32'h3f0cac9e : _GEN_595; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_5_io_in_b_Re = 5'h1a == _T_64[4:0] ? io_in_26_Re : _GEN_649; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_5_io_in_b_Im = 5'h1a == _T_64[4:0] ? io_in_26_Im : _GEN_622; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_io_in_a_Re = 5'h1a == _T_76[4:0] ? 32'hbf55e286 : _GEN_676; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_6_io_in_a_Im = 5'h1a == _T_76[4:0] ? 32'h3f0cac9e : _GEN_703; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_6_io_in_b_Re = 5'h1a == _T_76[4:0] ? io_in_26_Re : _GEN_757; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_6_io_in_b_Im = 5'h1a == _T_76[4:0] ? io_in_26_Im : _GEN_730; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_io_in_a_Re = 5'h1a == _T_88[4:0] ? 32'hbf55e286 : _GEN_784; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_7_io_in_a_Im = 5'h1a == _T_88[4:0] ? 32'h3f0cac9e : _GEN_811; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_7_io_in_b_Re = 5'h1a == _T_88[4:0] ? io_in_26_Re : _GEN_865; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_7_io_in_b_Im = 5'h1a == _T_88[4:0] ? io_in_26_Im : _GEN_838; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_io_in_a_Re = 5'h1a == _T_100[4:0] ? 32'hbf55e286 : _GEN_892; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_8_io_in_a_Im = 5'h1a == _T_100[4:0] ? 32'h3f0cac9e : _GEN_919; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_8_io_in_b_Re = 5'h1a == _T_100[4:0] ? io_in_26_Re : _GEN_973; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_8_io_in_b_Im = 5'h1a == _T_100[4:0] ? io_in_26_Im : _GEN_946; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_io_in_a_Re = 5'h1a == _T_112[4:0] ? 32'hbf55e286 : _GEN_1000; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_9_io_in_a_Im = 5'h1a == _T_112[4:0] ? 32'h3f0cac9e : _GEN_1027; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_9_io_in_b_Re = 5'h1a == _T_112[4:0] ? io_in_26_Re : _GEN_1081; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_9_io_in_b_Im = 5'h1a == _T_112[4:0] ? io_in_26_Im : _GEN_1054; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_io_in_a_Re = 5'h1a == _T_124[4:0] ? 32'hbf55e286 : _GEN_1108; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_10_io_in_a_Im = 5'h1a == _T_124[4:0] ? 32'h3f0cac9e : _GEN_1135; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_10_io_in_b_Re = 5'h1a == _T_124[4:0] ? io_in_26_Re : _GEN_1189; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_10_io_in_b_Im = 5'h1a == _T_124[4:0] ? io_in_26_Im : _GEN_1162; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_io_in_a_Re = 5'h1a == _T_136[4:0] ? 32'hbf55e286 : _GEN_1216; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_11_io_in_a_Im = 5'h1a == _T_136[4:0] ? 32'h3f0cac9e : _GEN_1243; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_11_io_in_b_Re = 5'h1a == _T_136[4:0] ? io_in_26_Re : _GEN_1297; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_11_io_in_b_Im = 5'h1a == _T_136[4:0] ? io_in_26_Im : _GEN_1270; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_12_clock = clock;
  assign FPComplexMult_12_io_in_a_Re = 5'h1a == _T_148[4:0] ? 32'hbf55e286 : _GEN_1324; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_12_io_in_a_Im = 5'h1a == _T_148[4:0] ? 32'h3f0cac9e : _GEN_1351; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_12_io_in_b_Re = 5'h1a == _T_148[4:0] ? io_in_26_Re : _GEN_1405; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_12_io_in_b_Im = 5'h1a == _T_148[4:0] ? io_in_26_Im : _GEN_1378; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_13_clock = clock;
  assign FPComplexMult_13_io_in_a_Re = 5'h1a == _T_160[4:0] ? 32'hbf55e286 : _GEN_1432; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_13_io_in_a_Im = 5'h1a == _T_160[4:0] ? 32'h3f0cac9e : _GEN_1459; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_13_io_in_b_Re = 5'h1a == _T_160[4:0] ? io_in_26_Re : _GEN_1513; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_13_io_in_b_Im = 5'h1a == _T_160[4:0] ? io_in_26_Im : _GEN_1486; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_14_clock = clock;
  assign FPComplexMult_14_io_in_a_Re = 5'h1a == _T_172[4:0] ? 32'hbf55e286 : _GEN_1540; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_14_io_in_a_Im = 5'h1a == _T_172[4:0] ? 32'h3f0cac9e : _GEN_1567; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_14_io_in_b_Re = 5'h1a == _T_172[4:0] ? io_in_26_Re : _GEN_1621; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_14_io_in_b_Im = 5'h1a == _T_172[4:0] ? io_in_26_Im : _GEN_1594; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_15_clock = clock;
  assign FPComplexMult_15_io_in_a_Re = 5'h1a == _T_184[4:0] ? 32'hbf55e286 : _GEN_1648; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_15_io_in_a_Im = 5'h1a == _T_184[4:0] ? 32'h3f0cac9e : _GEN_1675; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_15_io_in_b_Re = 5'h1a == _T_184[4:0] ? io_in_26_Re : _GEN_1729; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_15_io_in_b_Im = 5'h1a == _T_184[4:0] ? io_in_26_Im : _GEN_1702; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_16_clock = clock;
  assign FPComplexMult_16_io_in_a_Re = 5'h1a == _T_196[4:0] ? 32'hbf55e286 : _GEN_1756; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_16_io_in_a_Im = 5'h1a == _T_196[4:0] ? 32'h3f0cac9e : _GEN_1783; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_16_io_in_b_Re = 5'h1a == _T_196[4:0] ? io_in_26_Re : _GEN_1837; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_16_io_in_b_Im = 5'h1a == _T_196[4:0] ? io_in_26_Im : _GEN_1810; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_17_clock = clock;
  assign FPComplexMult_17_io_in_a_Re = 5'h1a == _T_208[4:0] ? 32'hbf55e286 : _GEN_1864; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_17_io_in_a_Im = 5'h1a == _T_208[4:0] ? 32'h3f0cac9e : _GEN_1891; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_17_io_in_b_Re = 5'h1a == _T_208[4:0] ? io_in_26_Re : _GEN_1945; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_17_io_in_b_Im = 5'h1a == _T_208[4:0] ? io_in_26_Im : _GEN_1918; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_18_clock = clock;
  assign FPComplexMult_18_io_in_a_Re = 5'h1a == _T_220[4:0] ? 32'hbf55e286 : _GEN_1972; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_18_io_in_a_Im = 5'h1a == _T_220[4:0] ? 32'h3f0cac9e : _GEN_1999; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_18_io_in_b_Re = 5'h1a == _T_220[4:0] ? io_in_26_Re : _GEN_2053; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_18_io_in_b_Im = 5'h1a == _T_220[4:0] ? io_in_26_Im : _GEN_2026; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_19_clock = clock;
  assign FPComplexMult_19_io_in_a_Re = 5'h1a == _T_232[4:0] ? 32'hbf55e286 : _GEN_2080; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_19_io_in_a_Im = 5'h1a == _T_232[4:0] ? 32'h3f0cac9e : _GEN_2107; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_19_io_in_b_Re = 5'h1a == _T_232[4:0] ? io_in_26_Re : _GEN_2161; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_19_io_in_b_Im = 5'h1a == _T_232[4:0] ? io_in_26_Im : _GEN_2134; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_20_clock = clock;
  assign FPComplexMult_20_io_in_a_Re = 5'h1a == _T_244[4:0] ? 32'hbf55e286 : _GEN_2188; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_20_io_in_a_Im = 5'h1a == _T_244[4:0] ? 32'h3f0cac9e : _GEN_2215; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_20_io_in_b_Re = 5'h1a == _T_244[4:0] ? io_in_26_Re : _GEN_2269; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_20_io_in_b_Im = 5'h1a == _T_244[4:0] ? io_in_26_Im : _GEN_2242; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_21_clock = clock;
  assign FPComplexMult_21_io_in_a_Re = 5'h1a == _T_256[4:0] ? 32'hbf55e286 : _GEN_2296; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_21_io_in_a_Im = 5'h1a == _T_256[4:0] ? 32'h3f0cac9e : _GEN_2323; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_21_io_in_b_Re = 5'h1a == _T_256[4:0] ? io_in_26_Re : _GEN_2377; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_21_io_in_b_Im = 5'h1a == _T_256[4:0] ? io_in_26_Im : _GEN_2350; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_22_clock = clock;
  assign FPComplexMult_22_io_in_a_Re = 5'h1a == _T_268[4:0] ? 32'hbf55e286 : _GEN_2404; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_22_io_in_a_Im = 5'h1a == _T_268[4:0] ? 32'h3f0cac9e : _GEN_2431; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_22_io_in_b_Re = 5'h1a == _T_268[4:0] ? io_in_26_Re : _GEN_2485; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_22_io_in_b_Im = 5'h1a == _T_268[4:0] ? io_in_26_Im : _GEN_2458; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_23_clock = clock;
  assign FPComplexMult_23_io_in_a_Re = 5'h1a == _T_280[4:0] ? 32'hbf55e286 : _GEN_2512; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_23_io_in_a_Im = 5'h1a == _T_280[4:0] ? 32'h3f0cac9e : _GEN_2539; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_23_io_in_b_Re = 5'h1a == _T_280[4:0] ? io_in_26_Re : _GEN_2593; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_23_io_in_b_Im = 5'h1a == _T_280[4:0] ? io_in_26_Im : _GEN_2566; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_24_clock = clock;
  assign FPComplexMult_24_io_in_a_Re = 5'h1a == _T_292[4:0] ? 32'hbf55e286 : _GEN_2620; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_24_io_in_a_Im = 5'h1a == _T_292[4:0] ? 32'h3f0cac9e : _GEN_2647; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_24_io_in_b_Re = 5'h1a == _T_292[4:0] ? io_in_26_Re : _GEN_2701; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_24_io_in_b_Im = 5'h1a == _T_292[4:0] ? io_in_26_Im : _GEN_2674; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_25_clock = clock;
  assign FPComplexMult_25_io_in_a_Re = 5'h1a == _T_304[4:0] ? 32'hbf55e286 : _GEN_2728; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_25_io_in_a_Im = 5'h1a == _T_304[4:0] ? 32'h3f0cac9e : _GEN_2755; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_25_io_in_b_Re = 5'h1a == _T_304[4:0] ? io_in_26_Re : _GEN_2809; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_25_io_in_b_Im = 5'h1a == _T_304[4:0] ? io_in_26_Im : _GEN_2782; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_26_clock = clock;
  assign FPComplexMult_26_io_in_a_Re = 5'h1a == _T_316[4:0] ? 32'hbf55e286 : _GEN_2836; // @[FFTDesigns.scala 541:{26,26}]
  assign FPComplexMult_26_io_in_a_Im = 5'h1a == _T_316[4:0] ? 32'h3f0cac9e : _GEN_2863; // @[FFTDesigns.scala 542:{26,26}]
  assign FPComplexMult_26_io_in_b_Re = 5'h1a == _T_316[4:0] ? io_in_26_Re : _GEN_2917; // @[FFTDesigns.scala 543:{23,23}]
  assign FPComplexMult_26_io_in_b_Im = 5'h1a == _T_316[4:0] ? io_in_26_Im : _GEN_2890; // @[FFTDesigns.scala 543:{23,23}]
  always @(posedge clock) begin
    if (cnt2 == 32'h1) begin // @[FFTDesigns.scala 529:38]
      if (cnt == 32'h0) begin // @[FFTDesigns.scala 531:32]
        cnt <= 32'h0; // @[FFTDesigns.scala 532:13]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 534:13]
      end
    end
    if (cnt2 == 32'h1) begin // @[FFTDesigns.scala 529:38]
      cnt2 <= 32'h0; // @[FFTDesigns.scala 530:12]
    end else begin
      cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 538:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cnt2 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FFT_sr(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input         io_in_ready,
  output        io_out_validate,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  DFT_r_V1_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_1_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_1_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_2_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_2_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_3_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_3_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_4_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_4_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_5_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_5_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_6_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_6_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_7_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_7_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_8_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_8_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_9_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_9_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_10_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_10_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_11_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_11_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_12_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_12_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_13_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_13_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_14_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_14_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_15_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_15_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_16_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_16_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_17_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_17_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_18_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_18_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_19_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_19_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_20_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_20_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_21_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_21_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_22_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_22_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_23_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_23_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_24_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_24_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_25_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_25_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire  DFT_r_V1_26_clock; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_in_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_in_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_in_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_in_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_in_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_in_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_out_0_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_out_0_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_out_1_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_out_1_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_out_2_Re; // @[FFTDesigns.scala 799:34]
  wire [31:0] DFT_r_V1_26_io_out_2_Im; // @[FFTDesigns.scala 799:34]
  wire [31:0] PermutationsBasic_io_in_0_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_0_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_1_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_1_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_2_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_2_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_3_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_3_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_4_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_4_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_5_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_5_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_6_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_6_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_7_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_7_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_8_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_8_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_9_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_9_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_10_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_10_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_11_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_11_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_12_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_12_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_13_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_13_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_14_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_14_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_15_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_15_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_16_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_16_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_17_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_17_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_18_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_18_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_19_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_19_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_20_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_20_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_21_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_21_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_22_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_22_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_23_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_23_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_24_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_24_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_25_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_25_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_26_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_in_26_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_3_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_3_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_4_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_4_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_5_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_5_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_6_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_6_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_7_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_7_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_8_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_8_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_9_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_9_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_10_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_10_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_11_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_11_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_12_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_12_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_13_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_13_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_14_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_14_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_15_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_15_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_16_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_16_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_17_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_17_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_18_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_18_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_19_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_19_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_20_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_20_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_21_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_21_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_22_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_22_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_23_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_23_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_24_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_24_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_25_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_25_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_26_Re; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_io_out_26_Im; // @[FFTDesigns.scala 804:35]
  wire [31:0] PermutationsBasic_1_io_in_0_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_0_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_1_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_1_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_2_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_2_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_3_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_3_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_4_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_4_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_5_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_5_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_6_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_6_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_7_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_7_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_8_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_8_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_9_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_9_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_10_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_10_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_11_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_11_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_12_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_12_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_13_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_13_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_14_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_14_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_15_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_15_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_16_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_16_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_17_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_17_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_18_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_18_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_19_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_19_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_20_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_20_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_21_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_21_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_22_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_22_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_23_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_23_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_24_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_24_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_25_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_25_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_26_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_in_26_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_3_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_3_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_4_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_4_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_5_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_5_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_6_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_6_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_7_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_7_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_8_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_8_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_9_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_9_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_10_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_10_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_11_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_11_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_12_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_12_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_13_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_13_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_14_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_14_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_15_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_15_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_16_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_16_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_17_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_17_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_18_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_18_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_19_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_19_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_20_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_20_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_21_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_21_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_22_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_22_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_23_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_23_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_24_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_24_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_25_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_25_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_26_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_1_io_out_26_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_0_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_0_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_1_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_1_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_2_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_2_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_3_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_3_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_4_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_4_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_5_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_5_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_6_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_6_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_7_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_7_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_8_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_8_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_9_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_9_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_10_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_10_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_11_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_11_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_12_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_12_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_13_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_13_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_14_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_14_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_15_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_15_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_16_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_16_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_17_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_17_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_18_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_18_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_19_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_19_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_20_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_20_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_21_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_21_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_22_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_22_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_23_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_23_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_24_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_24_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_25_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_25_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_26_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_in_26_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_0_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_0_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_1_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_1_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_2_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_2_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_3_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_3_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_4_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_4_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_5_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_5_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_6_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_6_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_7_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_7_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_8_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_8_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_9_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_9_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_10_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_10_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_11_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_11_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_12_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_12_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_13_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_13_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_14_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_14_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_15_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_15_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_16_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_16_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_17_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_17_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_18_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_18_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_19_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_19_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_20_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_20_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_21_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_21_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_22_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_22_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_23_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_23_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_24_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_24_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_25_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_25_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_26_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_2_io_out_26_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_0_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_0_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_1_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_1_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_2_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_2_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_3_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_3_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_4_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_4_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_5_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_5_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_6_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_6_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_7_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_7_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_8_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_8_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_9_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_9_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_10_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_10_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_11_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_11_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_12_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_12_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_13_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_13_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_14_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_14_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_15_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_15_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_16_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_16_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_17_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_17_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_18_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_18_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_19_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_19_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_20_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_20_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_21_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_21_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_22_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_22_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_23_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_23_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_24_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_24_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_25_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_25_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_26_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_in_26_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_0_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_0_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_1_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_1_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_2_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_2_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_3_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_3_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_4_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_4_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_5_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_5_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_6_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_6_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_7_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_7_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_8_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_8_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_9_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_9_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_10_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_10_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_11_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_11_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_12_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_12_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_13_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_13_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_14_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_14_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_15_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_15_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_16_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_16_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_17_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_17_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_18_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_18_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_19_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_19_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_20_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_20_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_21_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_21_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_22_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_22_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_23_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_23_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_24_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_24_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_25_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_25_Im; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_26_Re; // @[FFTDesigns.scala 806:37]
  wire [31:0] PermutationsBasic_3_io_out_26_Im; // @[FFTDesigns.scala 806:37]
  wire  TwiddleFactors_clock; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_0_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_0_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_1_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_1_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_2_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_2_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_3_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_3_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_4_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_4_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_5_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_5_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_6_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_6_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_7_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_7_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_8_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_8_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_9_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_9_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_10_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_10_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_11_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_11_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_12_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_12_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_13_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_13_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_14_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_14_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_15_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_15_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_16_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_16_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_17_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_17_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_18_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_18_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_19_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_19_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_20_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_20_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_21_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_21_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_22_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_22_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_23_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_23_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_24_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_24_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_25_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_25_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_26_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_in_26_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_0_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_0_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_1_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_1_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_2_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_2_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_3_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_3_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_4_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_4_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_5_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_5_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_6_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_6_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_7_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_7_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_8_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_8_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_9_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_9_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_10_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_10_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_11_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_11_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_12_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_12_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_13_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_13_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_14_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_14_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_15_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_15_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_16_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_16_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_17_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_17_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_18_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_18_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_19_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_19_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_20_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_20_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_21_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_21_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_22_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_22_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_23_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_23_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_24_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_24_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_25_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_25_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_26_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_io_out_26_Im; // @[FFTDesigns.scala 810:24]
  wire  TwiddleFactors_1_clock; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_0_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_0_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_1_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_1_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_2_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_2_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_3_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_3_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_4_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_4_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_5_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_5_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_6_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_6_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_7_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_7_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_8_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_8_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_9_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_9_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_10_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_10_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_11_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_11_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_12_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_12_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_13_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_13_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_14_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_14_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_15_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_15_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_16_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_16_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_17_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_17_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_18_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_18_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_19_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_19_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_20_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_20_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_21_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_21_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_22_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_22_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_23_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_23_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_24_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_24_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_25_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_25_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_26_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_in_26_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_0_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_0_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_1_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_1_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_2_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_2_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_3_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_3_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_4_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_4_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_5_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_5_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_6_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_6_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_7_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_7_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_8_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_8_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_9_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_9_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_10_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_10_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_11_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_11_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_12_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_12_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_13_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_13_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_14_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_14_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_15_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_15_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_16_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_16_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_17_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_17_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_18_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_18_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_19_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_19_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_20_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_20_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_21_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_21_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_22_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_22_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_23_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_23_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_24_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_24_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_25_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_25_Im; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_26_Re; // @[FFTDesigns.scala 810:24]
  wire [31:0] TwiddleFactors_1_io_out_26_Im; // @[FFTDesigns.scala 810:24]
  reg  regDelays_0; // @[FFTDesigns.scala 785:24]
  reg  regDelays_1; // @[FFTDesigns.scala 785:24]
  reg  regDelays_2; // @[FFTDesigns.scala 785:24]
  reg  regDelays_3; // @[FFTDesigns.scala 785:24]
  reg  regDelays_4; // @[FFTDesigns.scala 785:24]
  reg  regDelays_5; // @[FFTDesigns.scala 785:24]
  reg  regDelays_6; // @[FFTDesigns.scala 785:24]
  reg  regDelays_7; // @[FFTDesigns.scala 785:24]
  reg  regDelays_8; // @[FFTDesigns.scala 785:24]
  reg  regDelays_9; // @[FFTDesigns.scala 785:24]
  reg  regDelays_10; // @[FFTDesigns.scala 785:24]
  reg  regDelays_11; // @[FFTDesigns.scala 785:24]
  reg  regDelays_12; // @[FFTDesigns.scala 785:24]
  reg  regDelays_13; // @[FFTDesigns.scala 785:24]
  reg  regDelays_14; // @[FFTDesigns.scala 785:24]
  reg  regDelays_15; // @[FFTDesigns.scala 785:24]
  reg  regDelays_16; // @[FFTDesigns.scala 785:24]
  reg  regDelays_17; // @[FFTDesigns.scala 785:24]
  reg  regDelays_18; // @[FFTDesigns.scala 785:24]
  DFT_r_V1 DFT_r_V1 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_clock),
    .io_in_0_Re(DFT_r_V1_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_1 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_1_clock),
    .io_in_0_Re(DFT_r_V1_1_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_1_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_1_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_1_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_1_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_1_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_1_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_1_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_1_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_1_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_1_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_1_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_2 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_2_clock),
    .io_in_0_Re(DFT_r_V1_2_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_2_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_2_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_2_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_2_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_2_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_2_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_2_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_2_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_2_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_2_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_2_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_3 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_3_clock),
    .io_in_0_Re(DFT_r_V1_3_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_3_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_3_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_3_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_3_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_3_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_3_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_3_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_3_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_3_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_3_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_3_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_4 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_4_clock),
    .io_in_0_Re(DFT_r_V1_4_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_4_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_4_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_4_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_4_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_4_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_4_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_4_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_4_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_4_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_4_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_4_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_5 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_5_clock),
    .io_in_0_Re(DFT_r_V1_5_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_5_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_5_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_5_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_5_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_5_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_5_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_5_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_5_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_5_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_5_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_5_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_6 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_6_clock),
    .io_in_0_Re(DFT_r_V1_6_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_6_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_6_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_6_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_6_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_6_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_6_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_6_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_6_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_6_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_6_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_6_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_7 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_7_clock),
    .io_in_0_Re(DFT_r_V1_7_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_7_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_7_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_7_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_7_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_7_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_7_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_7_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_7_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_7_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_7_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_7_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_8 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_8_clock),
    .io_in_0_Re(DFT_r_V1_8_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_8_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_8_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_8_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_8_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_8_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_8_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_8_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_8_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_8_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_8_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_8_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_9 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_9_clock),
    .io_in_0_Re(DFT_r_V1_9_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_9_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_9_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_9_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_9_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_9_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_9_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_9_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_9_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_9_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_9_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_9_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_10 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_10_clock),
    .io_in_0_Re(DFT_r_V1_10_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_10_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_10_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_10_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_10_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_10_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_10_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_10_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_10_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_10_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_10_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_10_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_11 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_11_clock),
    .io_in_0_Re(DFT_r_V1_11_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_11_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_11_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_11_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_11_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_11_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_11_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_11_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_11_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_11_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_11_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_11_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_12 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_12_clock),
    .io_in_0_Re(DFT_r_V1_12_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_12_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_12_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_12_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_12_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_12_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_12_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_12_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_12_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_12_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_12_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_12_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_13 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_13_clock),
    .io_in_0_Re(DFT_r_V1_13_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_13_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_13_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_13_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_13_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_13_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_13_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_13_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_13_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_13_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_13_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_13_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_14 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_14_clock),
    .io_in_0_Re(DFT_r_V1_14_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_14_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_14_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_14_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_14_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_14_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_14_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_14_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_14_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_14_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_14_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_14_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_15 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_15_clock),
    .io_in_0_Re(DFT_r_V1_15_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_15_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_15_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_15_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_15_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_15_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_15_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_15_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_15_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_15_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_15_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_15_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_16 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_16_clock),
    .io_in_0_Re(DFT_r_V1_16_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_16_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_16_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_16_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_16_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_16_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_16_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_16_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_16_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_16_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_16_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_16_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_17 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_17_clock),
    .io_in_0_Re(DFT_r_V1_17_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_17_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_17_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_17_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_17_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_17_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_17_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_17_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_17_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_17_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_17_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_17_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_18 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_18_clock),
    .io_in_0_Re(DFT_r_V1_18_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_18_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_18_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_18_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_18_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_18_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_18_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_18_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_18_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_18_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_18_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_18_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_19 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_19_clock),
    .io_in_0_Re(DFT_r_V1_19_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_19_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_19_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_19_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_19_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_19_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_19_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_19_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_19_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_19_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_19_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_19_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_20 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_20_clock),
    .io_in_0_Re(DFT_r_V1_20_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_20_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_20_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_20_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_20_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_20_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_20_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_20_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_20_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_20_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_20_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_20_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_21 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_21_clock),
    .io_in_0_Re(DFT_r_V1_21_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_21_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_21_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_21_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_21_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_21_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_21_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_21_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_21_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_21_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_21_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_21_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_22 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_22_clock),
    .io_in_0_Re(DFT_r_V1_22_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_22_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_22_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_22_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_22_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_22_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_22_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_22_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_22_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_22_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_22_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_22_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_23 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_23_clock),
    .io_in_0_Re(DFT_r_V1_23_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_23_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_23_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_23_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_23_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_23_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_23_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_23_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_23_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_23_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_23_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_23_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_24 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_24_clock),
    .io_in_0_Re(DFT_r_V1_24_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_24_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_24_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_24_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_24_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_24_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_24_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_24_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_24_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_24_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_24_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_24_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_25 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_25_clock),
    .io_in_0_Re(DFT_r_V1_25_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_25_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_25_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_25_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_25_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_25_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_25_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_25_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_25_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_25_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_25_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_25_io_out_2_Im)
  );
  DFT_r_V1 DFT_r_V1_26 ( // @[FFTDesigns.scala 799:34]
    .clock(DFT_r_V1_26_clock),
    .io_in_0_Re(DFT_r_V1_26_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_26_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_26_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_26_io_in_1_Im),
    .io_in_2_Re(DFT_r_V1_26_io_in_2_Re),
    .io_in_2_Im(DFT_r_V1_26_io_in_2_Im),
    .io_out_0_Re(DFT_r_V1_26_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_26_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_26_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_26_io_out_1_Im),
    .io_out_2_Re(DFT_r_V1_26_io_out_2_Re),
    .io_out_2_Im(DFT_r_V1_26_io_out_2_Im)
  );
  PermutationsBasic PermutationsBasic ( // @[FFTDesigns.scala 804:35]
    .io_in_0_Re(PermutationsBasic_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_io_in_26_Im),
    .io_out_0_Re(PermutationsBasic_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_io_out_26_Im)
  );
  PermutationsBasic_1 PermutationsBasic_1 ( // @[FFTDesigns.scala 806:37]
    .io_in_0_Re(PermutationsBasic_1_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_1_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_1_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_1_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_1_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_1_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_1_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_1_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_1_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_1_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_1_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_1_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_1_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_1_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_1_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_1_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_1_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_1_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_1_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_1_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_1_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_1_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_1_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_1_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_1_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_1_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_1_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_1_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_1_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_1_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_1_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_1_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_1_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_1_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_1_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_1_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_1_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_1_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_1_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_1_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_1_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_1_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_1_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_1_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_1_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_1_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_1_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_1_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_1_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_1_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_1_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_1_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_1_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_1_io_in_26_Im),
    .io_out_0_Re(PermutationsBasic_1_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_1_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_1_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_1_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_1_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_1_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_1_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_1_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_1_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_1_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_1_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_1_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_1_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_1_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_1_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_1_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_1_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_1_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_1_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_1_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_1_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_1_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_1_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_1_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_1_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_1_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_1_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_1_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_1_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_1_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_1_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_1_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_1_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_1_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_1_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_1_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_1_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_1_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_1_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_1_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_1_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_1_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_1_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_1_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_1_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_1_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_1_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_1_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_1_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_1_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_1_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_1_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_1_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_1_io_out_26_Im)
  );
  PermutationsBasic_1 PermutationsBasic_2 ( // @[FFTDesigns.scala 806:37]
    .io_in_0_Re(PermutationsBasic_2_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_2_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_2_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_2_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_2_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_2_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_2_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_2_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_2_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_2_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_2_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_2_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_2_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_2_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_2_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_2_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_2_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_2_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_2_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_2_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_2_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_2_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_2_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_2_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_2_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_2_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_2_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_2_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_2_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_2_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_2_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_2_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_2_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_2_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_2_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_2_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_2_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_2_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_2_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_2_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_2_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_2_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_2_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_2_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_2_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_2_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_2_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_2_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_2_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_2_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_2_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_2_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_2_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_2_io_in_26_Im),
    .io_out_0_Re(PermutationsBasic_2_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_2_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_2_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_2_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_2_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_2_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_2_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_2_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_2_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_2_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_2_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_2_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_2_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_2_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_2_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_2_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_2_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_2_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_2_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_2_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_2_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_2_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_2_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_2_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_2_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_2_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_2_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_2_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_2_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_2_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_2_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_2_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_2_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_2_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_2_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_2_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_2_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_2_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_2_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_2_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_2_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_2_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_2_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_2_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_2_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_2_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_2_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_2_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_2_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_2_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_2_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_2_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_2_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_2_io_out_26_Im)
  );
  PermutationsBasic_1 PermutationsBasic_3 ( // @[FFTDesigns.scala 806:37]
    .io_in_0_Re(PermutationsBasic_3_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_3_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_3_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_3_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_3_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_3_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_3_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_3_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_3_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_3_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_3_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_3_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_3_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_3_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_3_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_3_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_3_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_3_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_3_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_3_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_3_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_3_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_3_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_3_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_3_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_3_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_3_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_3_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_3_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_3_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_3_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_3_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_3_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_3_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_3_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_3_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_3_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_3_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_3_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_3_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_3_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_3_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_3_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_3_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_3_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_3_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_3_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_3_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_3_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_3_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_3_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_3_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_3_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_3_io_in_26_Im),
    .io_out_0_Re(PermutationsBasic_3_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_3_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_3_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_3_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_3_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_3_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_3_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_3_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_3_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_3_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_3_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_3_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_3_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_3_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_3_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_3_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_3_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_3_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_3_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_3_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_3_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_3_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_3_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_3_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_3_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_3_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_3_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_3_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_3_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_3_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_3_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_3_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_3_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_3_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_3_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_3_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_3_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_3_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_3_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_3_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_3_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_3_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_3_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_3_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_3_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_3_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_3_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_3_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_3_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_3_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_3_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_3_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_3_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_3_io_out_26_Im)
  );
  TwiddleFactors TwiddleFactors ( // @[FFTDesigns.scala 810:24]
    .clock(TwiddleFactors_clock),
    .io_in_0_Re(TwiddleFactors_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_io_in_26_Im),
    .io_out_0_Re(TwiddleFactors_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_io_out_26_Im)
  );
  TwiddleFactors_1 TwiddleFactors_1 ( // @[FFTDesigns.scala 810:24]
    .clock(TwiddleFactors_1_clock),
    .io_in_0_Re(TwiddleFactors_1_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_1_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_1_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_1_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_1_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_1_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_1_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_1_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_1_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_1_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_1_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_1_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_1_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_1_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_1_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_1_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_1_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_1_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_1_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_1_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_1_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_1_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_1_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_1_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_1_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_1_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_1_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_1_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_1_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_1_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_1_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_1_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_1_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_1_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_1_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_1_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_1_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_1_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_1_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_1_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_1_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_1_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_1_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_1_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_1_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_1_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_1_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_1_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_1_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_1_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_1_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_1_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_1_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_1_io_in_26_Im),
    .io_out_0_Re(TwiddleFactors_1_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_1_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_1_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_1_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_1_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_1_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_1_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_1_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_1_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_1_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_1_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_1_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_1_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_1_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_1_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_1_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_1_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_1_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_1_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_1_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_1_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_1_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_1_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_1_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_1_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_1_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_1_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_1_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_1_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_1_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_1_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_1_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_1_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_1_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_1_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_1_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_1_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_1_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_1_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_1_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_1_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_1_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_1_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_1_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_1_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_1_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_1_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_1_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_1_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_1_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_1_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_1_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_1_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_1_io_out_26_Im)
  );
  assign io_out_validate = regDelays_18; // @[FFTDesigns.scala 793:28 794:18]
  assign io_out_0_Re = io_out_validate ? PermutationsBasic_3_io_out_0_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_0_Im = io_out_validate ? PermutationsBasic_3_io_out_0_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_1_Re = io_out_validate ? PermutationsBasic_3_io_out_1_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_1_Im = io_out_validate ? PermutationsBasic_3_io_out_1_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_2_Re = io_out_validate ? PermutationsBasic_3_io_out_2_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_2_Im = io_out_validate ? PermutationsBasic_3_io_out_2_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_3_Re = io_out_validate ? PermutationsBasic_3_io_out_3_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_3_Im = io_out_validate ? PermutationsBasic_3_io_out_3_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_4_Re = io_out_validate ? PermutationsBasic_3_io_out_4_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_4_Im = io_out_validate ? PermutationsBasic_3_io_out_4_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_5_Re = io_out_validate ? PermutationsBasic_3_io_out_5_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_5_Im = io_out_validate ? PermutationsBasic_3_io_out_5_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_6_Re = io_out_validate ? PermutationsBasic_3_io_out_6_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_6_Im = io_out_validate ? PermutationsBasic_3_io_out_6_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_7_Re = io_out_validate ? PermutationsBasic_3_io_out_7_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_7_Im = io_out_validate ? PermutationsBasic_3_io_out_7_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_8_Re = io_out_validate ? PermutationsBasic_3_io_out_8_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_8_Im = io_out_validate ? PermutationsBasic_3_io_out_8_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_9_Re = io_out_validate ? PermutationsBasic_3_io_out_9_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_9_Im = io_out_validate ? PermutationsBasic_3_io_out_9_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_10_Re = io_out_validate ? PermutationsBasic_3_io_out_10_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_10_Im = io_out_validate ? PermutationsBasic_3_io_out_10_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_11_Re = io_out_validate ? PermutationsBasic_3_io_out_11_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_11_Im = io_out_validate ? PermutationsBasic_3_io_out_11_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_12_Re = io_out_validate ? PermutationsBasic_3_io_out_12_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_12_Im = io_out_validate ? PermutationsBasic_3_io_out_12_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_13_Re = io_out_validate ? PermutationsBasic_3_io_out_13_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_13_Im = io_out_validate ? PermutationsBasic_3_io_out_13_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_14_Re = io_out_validate ? PermutationsBasic_3_io_out_14_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_14_Im = io_out_validate ? PermutationsBasic_3_io_out_14_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_15_Re = io_out_validate ? PermutationsBasic_3_io_out_15_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_15_Im = io_out_validate ? PermutationsBasic_3_io_out_15_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_16_Re = io_out_validate ? PermutationsBasic_3_io_out_16_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_16_Im = io_out_validate ? PermutationsBasic_3_io_out_16_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_17_Re = io_out_validate ? PermutationsBasic_3_io_out_17_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_17_Im = io_out_validate ? PermutationsBasic_3_io_out_17_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_18_Re = io_out_validate ? PermutationsBasic_3_io_out_18_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_18_Im = io_out_validate ? PermutationsBasic_3_io_out_18_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_19_Re = io_out_validate ? PermutationsBasic_3_io_out_19_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_19_Im = io_out_validate ? PermutationsBasic_3_io_out_19_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_20_Re = io_out_validate ? PermutationsBasic_3_io_out_20_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_20_Im = io_out_validate ? PermutationsBasic_3_io_out_20_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_21_Re = io_out_validate ? PermutationsBasic_3_io_out_21_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_21_Im = io_out_validate ? PermutationsBasic_3_io_out_21_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_22_Re = io_out_validate ? PermutationsBasic_3_io_out_22_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_22_Im = io_out_validate ? PermutationsBasic_3_io_out_22_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_23_Re = io_out_validate ? PermutationsBasic_3_io_out_23_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_23_Im = io_out_validate ? PermutationsBasic_3_io_out_23_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_24_Re = io_out_validate ? PermutationsBasic_3_io_out_24_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_24_Im = io_out_validate ? PermutationsBasic_3_io_out_24_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_25_Re = io_out_validate ? PermutationsBasic_3_io_out_25_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_25_Im = io_out_validate ? PermutationsBasic_3_io_out_25_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign io_out_26_Re = io_out_validate ? PermutationsBasic_3_io_out_26_Re : 32'h0; // @[FFTDesigns.scala 837:28 839:18 844:26]
  assign io_out_26_Im = io_out_validate ? PermutationsBasic_3_io_out_26_Im : 32'h0; // @[FFTDesigns.scala 837:28 839:18 845:26]
  assign DFT_r_V1_clock = clock;
  assign DFT_r_V1_io_in_0_Re = PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_io_in_0_Im = PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_io_in_1_Re = PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_io_in_1_Im = PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_io_in_2_Re = PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_io_in_2_Im = PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_1_clock = clock;
  assign DFT_r_V1_1_io_in_0_Re = PermutationsBasic_io_out_3_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_1_io_in_0_Im = PermutationsBasic_io_out_3_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_1_io_in_1_Re = PermutationsBasic_io_out_4_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_1_io_in_1_Im = PermutationsBasic_io_out_4_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_1_io_in_2_Re = PermutationsBasic_io_out_5_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_1_io_in_2_Im = PermutationsBasic_io_out_5_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_2_clock = clock;
  assign DFT_r_V1_2_io_in_0_Re = PermutationsBasic_io_out_6_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_2_io_in_0_Im = PermutationsBasic_io_out_6_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_2_io_in_1_Re = PermutationsBasic_io_out_7_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_2_io_in_1_Im = PermutationsBasic_io_out_7_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_2_io_in_2_Re = PermutationsBasic_io_out_8_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_2_io_in_2_Im = PermutationsBasic_io_out_8_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_3_clock = clock;
  assign DFT_r_V1_3_io_in_0_Re = PermutationsBasic_io_out_9_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_3_io_in_0_Im = PermutationsBasic_io_out_9_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_3_io_in_1_Re = PermutationsBasic_io_out_10_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_3_io_in_1_Im = PermutationsBasic_io_out_10_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_3_io_in_2_Re = PermutationsBasic_io_out_11_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_3_io_in_2_Im = PermutationsBasic_io_out_11_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_4_clock = clock;
  assign DFT_r_V1_4_io_in_0_Re = PermutationsBasic_io_out_12_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_4_io_in_0_Im = PermutationsBasic_io_out_12_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_4_io_in_1_Re = PermutationsBasic_io_out_13_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_4_io_in_1_Im = PermutationsBasic_io_out_13_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_4_io_in_2_Re = PermutationsBasic_io_out_14_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_4_io_in_2_Im = PermutationsBasic_io_out_14_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_5_clock = clock;
  assign DFT_r_V1_5_io_in_0_Re = PermutationsBasic_io_out_15_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_5_io_in_0_Im = PermutationsBasic_io_out_15_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_5_io_in_1_Re = PermutationsBasic_io_out_16_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_5_io_in_1_Im = PermutationsBasic_io_out_16_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_5_io_in_2_Re = PermutationsBasic_io_out_17_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_5_io_in_2_Im = PermutationsBasic_io_out_17_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_6_clock = clock;
  assign DFT_r_V1_6_io_in_0_Re = PermutationsBasic_io_out_18_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_6_io_in_0_Im = PermutationsBasic_io_out_18_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_6_io_in_1_Re = PermutationsBasic_io_out_19_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_6_io_in_1_Im = PermutationsBasic_io_out_19_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_6_io_in_2_Re = PermutationsBasic_io_out_20_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_6_io_in_2_Im = PermutationsBasic_io_out_20_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_7_clock = clock;
  assign DFT_r_V1_7_io_in_0_Re = PermutationsBasic_io_out_21_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_7_io_in_0_Im = PermutationsBasic_io_out_21_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_7_io_in_1_Re = PermutationsBasic_io_out_22_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_7_io_in_1_Im = PermutationsBasic_io_out_22_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_7_io_in_2_Re = PermutationsBasic_io_out_23_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_7_io_in_2_Im = PermutationsBasic_io_out_23_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_8_clock = clock;
  assign DFT_r_V1_8_io_in_0_Re = PermutationsBasic_io_out_24_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_8_io_in_0_Im = PermutationsBasic_io_out_24_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_8_io_in_1_Re = PermutationsBasic_io_out_25_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_8_io_in_1_Im = PermutationsBasic_io_out_25_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_8_io_in_2_Re = PermutationsBasic_io_out_26_Re; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_8_io_in_2_Im = PermutationsBasic_io_out_26_Im; // @[FFTDesigns.scala 827:39]
  assign DFT_r_V1_9_clock = clock;
  assign DFT_r_V1_9_io_in_0_Re = TwiddleFactors_io_out_0_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_9_io_in_0_Im = TwiddleFactors_io_out_0_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_9_io_in_1_Re = TwiddleFactors_io_out_1_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_9_io_in_1_Im = TwiddleFactors_io_out_1_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_9_io_in_2_Re = TwiddleFactors_io_out_2_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_9_io_in_2_Im = TwiddleFactors_io_out_2_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_10_clock = clock;
  assign DFT_r_V1_10_io_in_0_Re = TwiddleFactors_io_out_3_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_10_io_in_0_Im = TwiddleFactors_io_out_3_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_10_io_in_1_Re = TwiddleFactors_io_out_4_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_10_io_in_1_Im = TwiddleFactors_io_out_4_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_10_io_in_2_Re = TwiddleFactors_io_out_5_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_10_io_in_2_Im = TwiddleFactors_io_out_5_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_11_clock = clock;
  assign DFT_r_V1_11_io_in_0_Re = TwiddleFactors_io_out_6_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_11_io_in_0_Im = TwiddleFactors_io_out_6_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_11_io_in_1_Re = TwiddleFactors_io_out_7_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_11_io_in_1_Im = TwiddleFactors_io_out_7_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_11_io_in_2_Re = TwiddleFactors_io_out_8_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_11_io_in_2_Im = TwiddleFactors_io_out_8_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_12_clock = clock;
  assign DFT_r_V1_12_io_in_0_Re = TwiddleFactors_io_out_9_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_12_io_in_0_Im = TwiddleFactors_io_out_9_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_12_io_in_1_Re = TwiddleFactors_io_out_10_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_12_io_in_1_Im = TwiddleFactors_io_out_10_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_12_io_in_2_Re = TwiddleFactors_io_out_11_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_12_io_in_2_Im = TwiddleFactors_io_out_11_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_13_clock = clock;
  assign DFT_r_V1_13_io_in_0_Re = TwiddleFactors_io_out_12_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_13_io_in_0_Im = TwiddleFactors_io_out_12_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_13_io_in_1_Re = TwiddleFactors_io_out_13_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_13_io_in_1_Im = TwiddleFactors_io_out_13_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_13_io_in_2_Re = TwiddleFactors_io_out_14_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_13_io_in_2_Im = TwiddleFactors_io_out_14_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_14_clock = clock;
  assign DFT_r_V1_14_io_in_0_Re = TwiddleFactors_io_out_15_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_14_io_in_0_Im = TwiddleFactors_io_out_15_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_14_io_in_1_Re = TwiddleFactors_io_out_16_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_14_io_in_1_Im = TwiddleFactors_io_out_16_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_14_io_in_2_Re = TwiddleFactors_io_out_17_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_14_io_in_2_Im = TwiddleFactors_io_out_17_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_15_clock = clock;
  assign DFT_r_V1_15_io_in_0_Re = TwiddleFactors_io_out_18_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_15_io_in_0_Im = TwiddleFactors_io_out_18_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_15_io_in_1_Re = TwiddleFactors_io_out_19_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_15_io_in_1_Im = TwiddleFactors_io_out_19_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_15_io_in_2_Re = TwiddleFactors_io_out_20_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_15_io_in_2_Im = TwiddleFactors_io_out_20_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_16_clock = clock;
  assign DFT_r_V1_16_io_in_0_Re = TwiddleFactors_io_out_21_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_16_io_in_0_Im = TwiddleFactors_io_out_21_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_16_io_in_1_Re = TwiddleFactors_io_out_22_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_16_io_in_1_Im = TwiddleFactors_io_out_22_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_16_io_in_2_Re = TwiddleFactors_io_out_23_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_16_io_in_2_Im = TwiddleFactors_io_out_23_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_17_clock = clock;
  assign DFT_r_V1_17_io_in_0_Re = TwiddleFactors_io_out_24_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_17_io_in_0_Im = TwiddleFactors_io_out_24_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_17_io_in_1_Re = TwiddleFactors_io_out_25_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_17_io_in_1_Im = TwiddleFactors_io_out_25_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_17_io_in_2_Re = TwiddleFactors_io_out_26_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_17_io_in_2_Im = TwiddleFactors_io_out_26_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_18_clock = clock;
  assign DFT_r_V1_18_io_in_0_Re = TwiddleFactors_1_io_out_0_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_18_io_in_0_Im = TwiddleFactors_1_io_out_0_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_18_io_in_1_Re = TwiddleFactors_1_io_out_1_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_18_io_in_1_Im = TwiddleFactors_1_io_out_1_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_18_io_in_2_Re = TwiddleFactors_1_io_out_2_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_18_io_in_2_Im = TwiddleFactors_1_io_out_2_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_19_clock = clock;
  assign DFT_r_V1_19_io_in_0_Re = TwiddleFactors_1_io_out_3_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_19_io_in_0_Im = TwiddleFactors_1_io_out_3_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_19_io_in_1_Re = TwiddleFactors_1_io_out_4_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_19_io_in_1_Im = TwiddleFactors_1_io_out_4_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_19_io_in_2_Re = TwiddleFactors_1_io_out_5_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_19_io_in_2_Im = TwiddleFactors_1_io_out_5_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_20_clock = clock;
  assign DFT_r_V1_20_io_in_0_Re = TwiddleFactors_1_io_out_6_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_20_io_in_0_Im = TwiddleFactors_1_io_out_6_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_20_io_in_1_Re = TwiddleFactors_1_io_out_7_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_20_io_in_1_Im = TwiddleFactors_1_io_out_7_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_20_io_in_2_Re = TwiddleFactors_1_io_out_8_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_20_io_in_2_Im = TwiddleFactors_1_io_out_8_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_21_clock = clock;
  assign DFT_r_V1_21_io_in_0_Re = TwiddleFactors_1_io_out_9_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_21_io_in_0_Im = TwiddleFactors_1_io_out_9_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_21_io_in_1_Re = TwiddleFactors_1_io_out_10_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_21_io_in_1_Im = TwiddleFactors_1_io_out_10_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_21_io_in_2_Re = TwiddleFactors_1_io_out_11_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_21_io_in_2_Im = TwiddleFactors_1_io_out_11_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_22_clock = clock;
  assign DFT_r_V1_22_io_in_0_Re = TwiddleFactors_1_io_out_12_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_22_io_in_0_Im = TwiddleFactors_1_io_out_12_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_22_io_in_1_Re = TwiddleFactors_1_io_out_13_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_22_io_in_1_Im = TwiddleFactors_1_io_out_13_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_22_io_in_2_Re = TwiddleFactors_1_io_out_14_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_22_io_in_2_Im = TwiddleFactors_1_io_out_14_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_23_clock = clock;
  assign DFT_r_V1_23_io_in_0_Re = TwiddleFactors_1_io_out_15_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_23_io_in_0_Im = TwiddleFactors_1_io_out_15_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_23_io_in_1_Re = TwiddleFactors_1_io_out_16_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_23_io_in_1_Im = TwiddleFactors_1_io_out_16_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_23_io_in_2_Re = TwiddleFactors_1_io_out_17_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_23_io_in_2_Im = TwiddleFactors_1_io_out_17_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_24_clock = clock;
  assign DFT_r_V1_24_io_in_0_Re = TwiddleFactors_1_io_out_18_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_24_io_in_0_Im = TwiddleFactors_1_io_out_18_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_24_io_in_1_Re = TwiddleFactors_1_io_out_19_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_24_io_in_1_Im = TwiddleFactors_1_io_out_19_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_24_io_in_2_Re = TwiddleFactors_1_io_out_20_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_24_io_in_2_Im = TwiddleFactors_1_io_out_20_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_25_clock = clock;
  assign DFT_r_V1_25_io_in_0_Re = TwiddleFactors_1_io_out_21_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_25_io_in_0_Im = TwiddleFactors_1_io_out_21_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_25_io_in_1_Re = TwiddleFactors_1_io_out_22_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_25_io_in_1_Im = TwiddleFactors_1_io_out_22_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_25_io_in_2_Re = TwiddleFactors_1_io_out_23_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_25_io_in_2_Im = TwiddleFactors_1_io_out_23_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_26_clock = clock;
  assign DFT_r_V1_26_io_in_0_Re = TwiddleFactors_1_io_out_24_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_26_io_in_0_Im = TwiddleFactors_1_io_out_24_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_26_io_in_1_Re = TwiddleFactors_1_io_out_25_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_26_io_in_1_Im = TwiddleFactors_1_io_out_25_Im; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_26_io_in_2_Re = TwiddleFactors_1_io_out_26_Re; // @[FFTDesigns.scala 829:39]
  assign DFT_r_V1_26_io_in_2_Im = TwiddleFactors_1_io_out_26_Im; // @[FFTDesigns.scala 829:39]
  assign PermutationsBasic_io_in_0_Re = io_in_ready ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_0_Im = io_in_ready ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_1_Re = io_in_ready ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_1_Im = io_in_ready ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_2_Re = io_in_ready ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_2_Im = io_in_ready ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_3_Re = io_in_ready ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_3_Im = io_in_ready ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_4_Re = io_in_ready ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_4_Im = io_in_ready ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_5_Re = io_in_ready ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_5_Im = io_in_ready ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_6_Re = io_in_ready ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_6_Im = io_in_ready ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_7_Re = io_in_ready ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_7_Im = io_in_ready ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_8_Re = io_in_ready ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_8_Im = io_in_ready ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_9_Re = io_in_ready ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_9_Im = io_in_ready ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_10_Re = io_in_ready ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_10_Im = io_in_ready ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_11_Re = io_in_ready ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_11_Im = io_in_ready ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_12_Re = io_in_ready ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_12_Im = io_in_ready ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_13_Re = io_in_ready ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_13_Im = io_in_ready ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_14_Re = io_in_ready ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_14_Im = io_in_ready ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_15_Re = io_in_ready ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_15_Im = io_in_ready ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_16_Re = io_in_ready ? io_in_16_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_16_Im = io_in_ready ? io_in_16_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_17_Re = io_in_ready ? io_in_17_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_17_Im = io_in_ready ? io_in_17_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_18_Re = io_in_ready ? io_in_18_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_18_Im = io_in_ready ? io_in_18_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_19_Re = io_in_ready ? io_in_19_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_19_Im = io_in_ready ? io_in_19_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_20_Re = io_in_ready ? io_in_20_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_20_Im = io_in_ready ? io_in_20_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_21_Re = io_in_ready ? io_in_21_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_21_Im = io_in_ready ? io_in_21_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_22_Re = io_in_ready ? io_in_22_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_22_Im = io_in_ready ? io_in_22_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_23_Re = io_in_ready ? io_in_23_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_23_Im = io_in_ready ? io_in_23_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_24_Re = io_in_ready ? io_in_24_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_24_Im = io_in_ready ? io_in_24_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_25_Re = io_in_ready ? io_in_25_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_25_Im = io_in_ready ? io_in_25_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_io_in_26_Re = io_in_ready ? io_in_26_Re : 32'h0; // @[FFTDesigns.scala 813:22 815:33 819:36]
  assign PermutationsBasic_io_in_26_Im = io_in_ready ? io_in_26_Im : 32'h0; // @[FFTDesigns.scala 813:22 815:33 820:36]
  assign PermutationsBasic_1_io_in_0_Re = DFT_r_V1_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_0_Im = DFT_r_V1_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_1_Re = DFT_r_V1_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_1_Im = DFT_r_V1_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_2_Re = DFT_r_V1_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_2_Im = DFT_r_V1_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_3_Re = DFT_r_V1_1_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_3_Im = DFT_r_V1_1_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_4_Re = DFT_r_V1_1_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_4_Im = DFT_r_V1_1_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_5_Re = DFT_r_V1_1_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_5_Im = DFT_r_V1_1_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_6_Re = DFT_r_V1_2_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_6_Im = DFT_r_V1_2_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_7_Re = DFT_r_V1_2_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_7_Im = DFT_r_V1_2_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_8_Re = DFT_r_V1_2_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_8_Im = DFT_r_V1_2_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_9_Re = DFT_r_V1_3_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_9_Im = DFT_r_V1_3_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_10_Re = DFT_r_V1_3_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_10_Im = DFT_r_V1_3_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_11_Re = DFT_r_V1_3_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_11_Im = DFT_r_V1_3_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_12_Re = DFT_r_V1_4_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_12_Im = DFT_r_V1_4_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_13_Re = DFT_r_V1_4_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_13_Im = DFT_r_V1_4_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_14_Re = DFT_r_V1_4_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_14_Im = DFT_r_V1_4_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_15_Re = DFT_r_V1_5_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_15_Im = DFT_r_V1_5_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_16_Re = DFT_r_V1_5_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_16_Im = DFT_r_V1_5_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_17_Re = DFT_r_V1_5_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_17_Im = DFT_r_V1_5_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_18_Re = DFT_r_V1_6_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_18_Im = DFT_r_V1_6_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_19_Re = DFT_r_V1_6_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_19_Im = DFT_r_V1_6_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_20_Re = DFT_r_V1_6_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_20_Im = DFT_r_V1_6_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_21_Re = DFT_r_V1_7_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_21_Im = DFT_r_V1_7_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_22_Re = DFT_r_V1_7_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_22_Im = DFT_r_V1_7_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_23_Re = DFT_r_V1_7_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_23_Im = DFT_r_V1_7_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_24_Re = DFT_r_V1_8_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_24_Im = DFT_r_V1_8_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_25_Re = DFT_r_V1_8_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_25_Im = DFT_r_V1_8_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_26_Re = DFT_r_V1_8_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_1_io_in_26_Im = DFT_r_V1_8_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_0_Re = DFT_r_V1_9_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_0_Im = DFT_r_V1_9_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_1_Re = DFT_r_V1_9_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_1_Im = DFT_r_V1_9_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_2_Re = DFT_r_V1_9_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_2_Im = DFT_r_V1_9_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_3_Re = DFT_r_V1_10_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_3_Im = DFT_r_V1_10_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_4_Re = DFT_r_V1_10_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_4_Im = DFT_r_V1_10_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_5_Re = DFT_r_V1_10_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_5_Im = DFT_r_V1_10_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_6_Re = DFT_r_V1_11_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_6_Im = DFT_r_V1_11_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_7_Re = DFT_r_V1_11_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_7_Im = DFT_r_V1_11_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_8_Re = DFT_r_V1_11_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_8_Im = DFT_r_V1_11_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_9_Re = DFT_r_V1_12_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_9_Im = DFT_r_V1_12_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_10_Re = DFT_r_V1_12_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_10_Im = DFT_r_V1_12_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_11_Re = DFT_r_V1_12_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_11_Im = DFT_r_V1_12_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_12_Re = DFT_r_V1_13_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_12_Im = DFT_r_V1_13_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_13_Re = DFT_r_V1_13_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_13_Im = DFT_r_V1_13_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_14_Re = DFT_r_V1_13_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_14_Im = DFT_r_V1_13_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_15_Re = DFT_r_V1_14_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_15_Im = DFT_r_V1_14_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_16_Re = DFT_r_V1_14_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_16_Im = DFT_r_V1_14_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_17_Re = DFT_r_V1_14_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_17_Im = DFT_r_V1_14_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_18_Re = DFT_r_V1_15_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_18_Im = DFT_r_V1_15_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_19_Re = DFT_r_V1_15_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_19_Im = DFT_r_V1_15_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_20_Re = DFT_r_V1_15_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_20_Im = DFT_r_V1_15_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_21_Re = DFT_r_V1_16_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_21_Im = DFT_r_V1_16_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_22_Re = DFT_r_V1_16_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_22_Im = DFT_r_V1_16_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_23_Re = DFT_r_V1_16_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_23_Im = DFT_r_V1_16_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_24_Re = DFT_r_V1_17_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_24_Im = DFT_r_V1_17_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_25_Re = DFT_r_V1_17_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_25_Im = DFT_r_V1_17_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_26_Re = DFT_r_V1_17_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_2_io_in_26_Im = DFT_r_V1_17_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_0_Re = DFT_r_V1_18_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_0_Im = DFT_r_V1_18_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_1_Re = DFT_r_V1_18_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_1_Im = DFT_r_V1_18_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_2_Re = DFT_r_V1_18_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_2_Im = DFT_r_V1_18_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_3_Re = DFT_r_V1_19_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_3_Im = DFT_r_V1_19_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_4_Re = DFT_r_V1_19_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_4_Im = DFT_r_V1_19_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_5_Re = DFT_r_V1_19_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_5_Im = DFT_r_V1_19_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_6_Re = DFT_r_V1_20_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_6_Im = DFT_r_V1_20_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_7_Re = DFT_r_V1_20_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_7_Im = DFT_r_V1_20_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_8_Re = DFT_r_V1_20_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_8_Im = DFT_r_V1_20_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_9_Re = DFT_r_V1_21_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_9_Im = DFT_r_V1_21_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_10_Re = DFT_r_V1_21_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_10_Im = DFT_r_V1_21_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_11_Re = DFT_r_V1_21_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_11_Im = DFT_r_V1_21_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_12_Re = DFT_r_V1_22_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_12_Im = DFT_r_V1_22_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_13_Re = DFT_r_V1_22_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_13_Im = DFT_r_V1_22_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_14_Re = DFT_r_V1_22_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_14_Im = DFT_r_V1_22_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_15_Re = DFT_r_V1_23_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_15_Im = DFT_r_V1_23_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_16_Re = DFT_r_V1_23_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_16_Im = DFT_r_V1_23_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_17_Re = DFT_r_V1_23_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_17_Im = DFT_r_V1_23_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_18_Re = DFT_r_V1_24_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_18_Im = DFT_r_V1_24_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_19_Re = DFT_r_V1_24_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_19_Im = DFT_r_V1_24_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_20_Re = DFT_r_V1_24_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_20_Im = DFT_r_V1_24_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_21_Re = DFT_r_V1_25_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_21_Im = DFT_r_V1_25_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_22_Re = DFT_r_V1_25_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_22_Im = DFT_r_V1_25_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_23_Re = DFT_r_V1_25_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_23_Im = DFT_r_V1_25_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_24_Re = DFT_r_V1_26_io_out_0_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_24_Im = DFT_r_V1_26_io_out_0_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_25_Re = DFT_r_V1_26_io_out_1_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_25_Im = DFT_r_V1_26_io_out_1_Im; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_26_Re = DFT_r_V1_26_io_out_2_Re; // @[FFTDesigns.scala 831:43]
  assign PermutationsBasic_3_io_in_26_Im = DFT_r_V1_26_io_out_2_Im; // @[FFTDesigns.scala 831:43]
  assign TwiddleFactors_clock = clock;
  assign TwiddleFactors_io_in_0_Re = PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_0_Im = PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_1_Re = PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_1_Im = PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_2_Re = PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_2_Im = PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_3_Re = PermutationsBasic_1_io_out_3_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_3_Im = PermutationsBasic_1_io_out_3_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_4_Re = PermutationsBasic_1_io_out_4_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_4_Im = PermutationsBasic_1_io_out_4_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_5_Re = PermutationsBasic_1_io_out_5_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_5_Im = PermutationsBasic_1_io_out_5_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_6_Re = PermutationsBasic_1_io_out_6_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_6_Im = PermutationsBasic_1_io_out_6_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_7_Re = PermutationsBasic_1_io_out_7_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_7_Im = PermutationsBasic_1_io_out_7_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_8_Re = PermutationsBasic_1_io_out_8_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_8_Im = PermutationsBasic_1_io_out_8_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_9_Re = PermutationsBasic_1_io_out_9_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_9_Im = PermutationsBasic_1_io_out_9_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_10_Re = PermutationsBasic_1_io_out_10_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_10_Im = PermutationsBasic_1_io_out_10_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_11_Re = PermutationsBasic_1_io_out_11_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_11_Im = PermutationsBasic_1_io_out_11_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_12_Re = PermutationsBasic_1_io_out_12_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_12_Im = PermutationsBasic_1_io_out_12_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_13_Re = PermutationsBasic_1_io_out_13_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_13_Im = PermutationsBasic_1_io_out_13_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_14_Re = PermutationsBasic_1_io_out_14_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_14_Im = PermutationsBasic_1_io_out_14_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_15_Re = PermutationsBasic_1_io_out_15_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_15_Im = PermutationsBasic_1_io_out_15_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_16_Re = PermutationsBasic_1_io_out_16_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_16_Im = PermutationsBasic_1_io_out_16_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_17_Re = PermutationsBasic_1_io_out_17_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_17_Im = PermutationsBasic_1_io_out_17_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_18_Re = PermutationsBasic_1_io_out_18_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_18_Im = PermutationsBasic_1_io_out_18_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_19_Re = PermutationsBasic_1_io_out_19_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_19_Im = PermutationsBasic_1_io_out_19_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_20_Re = PermutationsBasic_1_io_out_20_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_20_Im = PermutationsBasic_1_io_out_20_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_21_Re = PermutationsBasic_1_io_out_21_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_21_Im = PermutationsBasic_1_io_out_21_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_22_Re = PermutationsBasic_1_io_out_22_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_22_Im = PermutationsBasic_1_io_out_22_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_23_Re = PermutationsBasic_1_io_out_23_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_23_Im = PermutationsBasic_1_io_out_23_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_24_Re = PermutationsBasic_1_io_out_24_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_24_Im = PermutationsBasic_1_io_out_24_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_25_Re = PermutationsBasic_1_io_out_25_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_25_Im = PermutationsBasic_1_io_out_25_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_26_Re = PermutationsBasic_1_io_out_26_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_io_in_26_Im = PermutationsBasic_1_io_out_26_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_clock = clock;
  assign TwiddleFactors_1_io_in_0_Re = PermutationsBasic_2_io_out_0_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_0_Im = PermutationsBasic_2_io_out_0_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_1_Re = PermutationsBasic_2_io_out_1_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_1_Im = PermutationsBasic_2_io_out_1_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_2_Re = PermutationsBasic_2_io_out_2_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_2_Im = PermutationsBasic_2_io_out_2_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_3_Re = PermutationsBasic_2_io_out_3_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_3_Im = PermutationsBasic_2_io_out_3_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_4_Re = PermutationsBasic_2_io_out_4_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_4_Im = PermutationsBasic_2_io_out_4_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_5_Re = PermutationsBasic_2_io_out_5_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_5_Im = PermutationsBasic_2_io_out_5_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_6_Re = PermutationsBasic_2_io_out_6_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_6_Im = PermutationsBasic_2_io_out_6_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_7_Re = PermutationsBasic_2_io_out_7_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_7_Im = PermutationsBasic_2_io_out_7_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_8_Re = PermutationsBasic_2_io_out_8_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_8_Im = PermutationsBasic_2_io_out_8_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_9_Re = PermutationsBasic_2_io_out_9_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_9_Im = PermutationsBasic_2_io_out_9_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_10_Re = PermutationsBasic_2_io_out_10_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_10_Im = PermutationsBasic_2_io_out_10_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_11_Re = PermutationsBasic_2_io_out_11_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_11_Im = PermutationsBasic_2_io_out_11_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_12_Re = PermutationsBasic_2_io_out_12_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_12_Im = PermutationsBasic_2_io_out_12_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_13_Re = PermutationsBasic_2_io_out_13_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_13_Im = PermutationsBasic_2_io_out_13_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_14_Re = PermutationsBasic_2_io_out_14_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_14_Im = PermutationsBasic_2_io_out_14_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_15_Re = PermutationsBasic_2_io_out_15_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_15_Im = PermutationsBasic_2_io_out_15_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_16_Re = PermutationsBasic_2_io_out_16_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_16_Im = PermutationsBasic_2_io_out_16_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_17_Re = PermutationsBasic_2_io_out_17_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_17_Im = PermutationsBasic_2_io_out_17_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_18_Re = PermutationsBasic_2_io_out_18_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_18_Im = PermutationsBasic_2_io_out_18_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_19_Re = PermutationsBasic_2_io_out_19_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_19_Im = PermutationsBasic_2_io_out_19_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_20_Re = PermutationsBasic_2_io_out_20_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_20_Im = PermutationsBasic_2_io_out_20_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_21_Re = PermutationsBasic_2_io_out_21_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_21_Im = PermutationsBasic_2_io_out_21_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_22_Re = PermutationsBasic_2_io_out_22_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_22_Im = PermutationsBasic_2_io_out_22_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_23_Re = PermutationsBasic_2_io_out_23_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_23_Im = PermutationsBasic_2_io_out_23_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_24_Re = PermutationsBasic_2_io_out_24_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_24_Im = PermutationsBasic_2_io_out_24_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_25_Re = PermutationsBasic_2_io_out_25_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_25_Im = PermutationsBasic_2_io_out_25_Im; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_26_Re = PermutationsBasic_2_io_out_26_Re; // @[FFTDesigns.scala 835:38]
  assign TwiddleFactors_1_io_in_26_Im = PermutationsBasic_2_io_out_26_Im; // @[FFTDesigns.scala 835:38]
  always @(posedge clock) begin
    regDelays_0 <= io_in_ready; // @[FFTDesigns.scala 788:22]
    regDelays_1 <= regDelays_0; // @[FFTDesigns.scala 790:22]
    regDelays_2 <= regDelays_1; // @[FFTDesigns.scala 790:22]
    regDelays_3 <= regDelays_2; // @[FFTDesigns.scala 790:22]
    regDelays_4 <= regDelays_3; // @[FFTDesigns.scala 790:22]
    regDelays_5 <= regDelays_4; // @[FFTDesigns.scala 790:22]
    regDelays_6 <= regDelays_5; // @[FFTDesigns.scala 790:22]
    regDelays_7 <= regDelays_6; // @[FFTDesigns.scala 790:22]
    regDelays_8 <= regDelays_7; // @[FFTDesigns.scala 790:22]
    regDelays_9 <= regDelays_8; // @[FFTDesigns.scala 790:22]
    regDelays_10 <= regDelays_9; // @[FFTDesigns.scala 790:22]
    regDelays_11 <= regDelays_10; // @[FFTDesigns.scala 790:22]
    regDelays_12 <= regDelays_11; // @[FFTDesigns.scala 790:22]
    regDelays_13 <= regDelays_12; // @[FFTDesigns.scala 790:22]
    regDelays_14 <= regDelays_13; // @[FFTDesigns.scala 790:22]
    regDelays_15 <= regDelays_14; // @[FFTDesigns.scala 790:22]
    regDelays_16 <= regDelays_15; // @[FFTDesigns.scala 790:22]
    regDelays_17 <= regDelays_16; // @[FFTDesigns.scala 790:22]
    regDelays_18 <= regDelays_17; // @[FFTDesigns.scala 790:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regDelays_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  regDelays_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  regDelays_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  regDelays_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  regDelays_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regDelays_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  regDelays_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  regDelays_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  regDelays_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  regDelays_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  regDelays_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  regDelays_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  regDelays_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  regDelays_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  regDelays_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  regDelays_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  regDelays_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  regDelays_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  regDelays_18 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

